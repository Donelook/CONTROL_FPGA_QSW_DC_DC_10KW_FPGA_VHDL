// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 12 2024 23:00:57

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    test,
    start_stop,
    s2_phy,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    clock_output,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    test22,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output test;
    input start_stop;
    output s2_phy;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output clock_output;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    output test22;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__51011;
    wire N__51010;
    wire N__51009;
    wire N__51000;
    wire N__50999;
    wire N__50998;
    wire N__50991;
    wire N__50990;
    wire N__50989;
    wire N__50982;
    wire N__50981;
    wire N__50980;
    wire N__50973;
    wire N__50972;
    wire N__50971;
    wire N__50964;
    wire N__50963;
    wire N__50962;
    wire N__50955;
    wire N__50954;
    wire N__50953;
    wire N__50946;
    wire N__50945;
    wire N__50944;
    wire N__50937;
    wire N__50936;
    wire N__50935;
    wire N__50928;
    wire N__50927;
    wire N__50926;
    wire N__50919;
    wire N__50918;
    wire N__50917;
    wire N__50910;
    wire N__50909;
    wire N__50908;
    wire N__50901;
    wire N__50900;
    wire N__50899;
    wire N__50892;
    wire N__50891;
    wire N__50890;
    wire N__50883;
    wire N__50882;
    wire N__50881;
    wire N__50874;
    wire N__50873;
    wire N__50872;
    wire N__50855;
    wire N__50852;
    wire N__50851;
    wire N__50850;
    wire N__50847;
    wire N__50844;
    wire N__50841;
    wire N__50836;
    wire N__50831;
    wire N__50828;
    wire N__50827;
    wire N__50824;
    wire N__50821;
    wire N__50820;
    wire N__50815;
    wire N__50812;
    wire N__50809;
    wire N__50804;
    wire N__50801;
    wire N__50800;
    wire N__50797;
    wire N__50794;
    wire N__50791;
    wire N__50786;
    wire N__50783;
    wire N__50782;
    wire N__50781;
    wire N__50780;
    wire N__50779;
    wire N__50778;
    wire N__50777;
    wire N__50776;
    wire N__50775;
    wire N__50774;
    wire N__50773;
    wire N__50772;
    wire N__50771;
    wire N__50770;
    wire N__50769;
    wire N__50768;
    wire N__50767;
    wire N__50766;
    wire N__50765;
    wire N__50764;
    wire N__50763;
    wire N__50762;
    wire N__50761;
    wire N__50760;
    wire N__50759;
    wire N__50758;
    wire N__50757;
    wire N__50756;
    wire N__50755;
    wire N__50754;
    wire N__50745;
    wire N__50736;
    wire N__50731;
    wire N__50722;
    wire N__50713;
    wire N__50704;
    wire N__50695;
    wire N__50686;
    wire N__50673;
    wire N__50668;
    wire N__50665;
    wire N__50660;
    wire N__50657;
    wire N__50656;
    wire N__50653;
    wire N__50650;
    wire N__50647;
    wire N__50642;
    wire N__50641;
    wire N__50640;
    wire N__50637;
    wire N__50634;
    wire N__50633;
    wire N__50630;
    wire N__50625;
    wire N__50622;
    wire N__50619;
    wire N__50616;
    wire N__50613;
    wire N__50610;
    wire N__50607;
    wire N__50604;
    wire N__50597;
    wire N__50594;
    wire N__50591;
    wire N__50590;
    wire N__50589;
    wire N__50588;
    wire N__50585;
    wire N__50580;
    wire N__50577;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50563;
    wire N__50558;
    wire N__50557;
    wire N__50556;
    wire N__50553;
    wire N__50550;
    wire N__50547;
    wire N__50544;
    wire N__50541;
    wire N__50536;
    wire N__50533;
    wire N__50528;
    wire N__50527;
    wire N__50526;
    wire N__50525;
    wire N__50524;
    wire N__50523;
    wire N__50522;
    wire N__50521;
    wire N__50520;
    wire N__50519;
    wire N__50518;
    wire N__50517;
    wire N__50516;
    wire N__50515;
    wire N__50514;
    wire N__50513;
    wire N__50512;
    wire N__50511;
    wire N__50510;
    wire N__50509;
    wire N__50508;
    wire N__50507;
    wire N__50506;
    wire N__50505;
    wire N__50502;
    wire N__50501;
    wire N__50500;
    wire N__50499;
    wire N__50498;
    wire N__50497;
    wire N__50496;
    wire N__50495;
    wire N__50494;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50486;
    wire N__50485;
    wire N__50484;
    wire N__50483;
    wire N__50482;
    wire N__50481;
    wire N__50480;
    wire N__50479;
    wire N__50478;
    wire N__50477;
    wire N__50474;
    wire N__50473;
    wire N__50470;
    wire N__50469;
    wire N__50464;
    wire N__50461;
    wire N__50458;
    wire N__50449;
    wire N__50442;
    wire N__50435;
    wire N__50424;
    wire N__50421;
    wire N__50420;
    wire N__50417;
    wire N__50412;
    wire N__50411;
    wire N__50410;
    wire N__50409;
    wire N__50408;
    wire N__50407;
    wire N__50406;
    wire N__50405;
    wire N__50404;
    wire N__50403;
    wire N__50402;
    wire N__50401;
    wire N__50400;
    wire N__50399;
    wire N__50398;
    wire N__50397;
    wire N__50396;
    wire N__50395;
    wire N__50394;
    wire N__50391;
    wire N__50390;
    wire N__50381;
    wire N__50378;
    wire N__50375;
    wire N__50372;
    wire N__50367;
    wire N__50364;
    wire N__50355;
    wire N__50354;
    wire N__50353;
    wire N__50352;
    wire N__50351;
    wire N__50340;
    wire N__50337;
    wire N__50334;
    wire N__50333;
    wire N__50332;
    wire N__50331;
    wire N__50330;
    wire N__50329;
    wire N__50328;
    wire N__50327;
    wire N__50326;
    wire N__50325;
    wire N__50322;
    wire N__50319;
    wire N__50314;
    wire N__50311;
    wire N__50304;
    wire N__50303;
    wire N__50302;
    wire N__50299;
    wire N__50298;
    wire N__50297;
    wire N__50296;
    wire N__50295;
    wire N__50294;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50283;
    wire N__50282;
    wire N__50281;
    wire N__50276;
    wire N__50265;
    wire N__50256;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50234;
    wire N__50219;
    wire N__50210;
    wire N__50207;
    wire N__50202;
    wire N__50189;
    wire N__50182;
    wire N__50173;
    wire N__50170;
    wire N__50165;
    wire N__50160;
    wire N__50151;
    wire N__50142;
    wire N__50137;
    wire N__50130;
    wire N__50123;
    wire N__50116;
    wire N__50111;
    wire N__50104;
    wire N__50075;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50063;
    wire N__50060;
    wire N__50057;
    wire N__50054;
    wire N__50051;
    wire N__50050;
    wire N__50049;
    wire N__50048;
    wire N__50047;
    wire N__50046;
    wire N__50045;
    wire N__50044;
    wire N__50043;
    wire N__50042;
    wire N__50041;
    wire N__50040;
    wire N__50039;
    wire N__50038;
    wire N__50037;
    wire N__50036;
    wire N__50035;
    wire N__50034;
    wire N__50033;
    wire N__50032;
    wire N__50031;
    wire N__50030;
    wire N__50029;
    wire N__50028;
    wire N__50027;
    wire N__50026;
    wire N__50025;
    wire N__50024;
    wire N__50023;
    wire N__50022;
    wire N__50021;
    wire N__50020;
    wire N__50019;
    wire N__50018;
    wire N__50017;
    wire N__50016;
    wire N__50015;
    wire N__50014;
    wire N__50013;
    wire N__50012;
    wire N__50011;
    wire N__50010;
    wire N__50009;
    wire N__50008;
    wire N__50007;
    wire N__50006;
    wire N__50005;
    wire N__50004;
    wire N__50003;
    wire N__50002;
    wire N__50001;
    wire N__50000;
    wire N__49999;
    wire N__49998;
    wire N__49997;
    wire N__49996;
    wire N__49995;
    wire N__49994;
    wire N__49993;
    wire N__49992;
    wire N__49991;
    wire N__49990;
    wire N__49989;
    wire N__49988;
    wire N__49987;
    wire N__49986;
    wire N__49985;
    wire N__49984;
    wire N__49983;
    wire N__49982;
    wire N__49981;
    wire N__49980;
    wire N__49979;
    wire N__49978;
    wire N__49977;
    wire N__49976;
    wire N__49975;
    wire N__49974;
    wire N__49973;
    wire N__49972;
    wire N__49971;
    wire N__49970;
    wire N__49969;
    wire N__49968;
    wire N__49967;
    wire N__49966;
    wire N__49965;
    wire N__49964;
    wire N__49963;
    wire N__49962;
    wire N__49961;
    wire N__49960;
    wire N__49959;
    wire N__49958;
    wire N__49957;
    wire N__49956;
    wire N__49955;
    wire N__49954;
    wire N__49953;
    wire N__49952;
    wire N__49951;
    wire N__49950;
    wire N__49949;
    wire N__49948;
    wire N__49947;
    wire N__49946;
    wire N__49945;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49941;
    wire N__49940;
    wire N__49939;
    wire N__49938;
    wire N__49937;
    wire N__49936;
    wire N__49935;
    wire N__49934;
    wire N__49933;
    wire N__49932;
    wire N__49931;
    wire N__49930;
    wire N__49929;
    wire N__49928;
    wire N__49927;
    wire N__49926;
    wire N__49925;
    wire N__49924;
    wire N__49923;
    wire N__49922;
    wire N__49921;
    wire N__49920;
    wire N__49919;
    wire N__49918;
    wire N__49917;
    wire N__49916;
    wire N__49915;
    wire N__49914;
    wire N__49913;
    wire N__49912;
    wire N__49911;
    wire N__49910;
    wire N__49909;
    wire N__49908;
    wire N__49907;
    wire N__49906;
    wire N__49905;
    wire N__49904;
    wire N__49903;
    wire N__49902;
    wire N__49901;
    wire N__49900;
    wire N__49899;
    wire N__49896;
    wire N__49895;
    wire N__49894;
    wire N__49583;
    wire N__49580;
    wire N__49579;
    wire N__49578;
    wire N__49577;
    wire N__49570;
    wire N__49567;
    wire N__49566;
    wire N__49565;
    wire N__49564;
    wire N__49563;
    wire N__49560;
    wire N__49557;
    wire N__49554;
    wire N__49551;
    wire N__49550;
    wire N__49549;
    wire N__49548;
    wire N__49545;
    wire N__49544;
    wire N__49543;
    wire N__49542;
    wire N__49539;
    wire N__49530;
    wire N__49529;
    wire N__49528;
    wire N__49527;
    wire N__49526;
    wire N__49525;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49521;
    wire N__49520;
    wire N__49517;
    wire N__49514;
    wire N__49511;
    wire N__49508;
    wire N__49505;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49497;
    wire N__49494;
    wire N__49491;
    wire N__49482;
    wire N__49473;
    wire N__49472;
    wire N__49471;
    wire N__49470;
    wire N__49469;
    wire N__49466;
    wire N__49465;
    wire N__49464;
    wire N__49463;
    wire N__49462;
    wire N__49461;
    wire N__49460;
    wire N__49457;
    wire N__49454;
    wire N__49451;
    wire N__49448;
    wire N__49443;
    wire N__49440;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49430;
    wire N__49429;
    wire N__49426;
    wire N__49417;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49393;
    wire N__49390;
    wire N__49389;
    wire N__49388;
    wire N__49387;
    wire N__49378;
    wire N__49375;
    wire N__49372;
    wire N__49369;
    wire N__49360;
    wire N__49359;
    wire N__49358;
    wire N__49357;
    wire N__49356;
    wire N__49353;
    wire N__49350;
    wire N__49347;
    wire N__49342;
    wire N__49339;
    wire N__49334;
    wire N__49331;
    wire N__49324;
    wire N__49321;
    wire N__49316;
    wire N__49311;
    wire N__49302;
    wire N__49297;
    wire N__49288;
    wire N__49271;
    wire N__49270;
    wire N__49269;
    wire N__49268;
    wire N__49265;
    wire N__49262;
    wire N__49259;
    wire N__49256;
    wire N__49253;
    wire N__49250;
    wire N__49247;
    wire N__49246;
    wire N__49245;
    wire N__49244;
    wire N__49241;
    wire N__49240;
    wire N__49239;
    wire N__49238;
    wire N__49237;
    wire N__49236;
    wire N__49235;
    wire N__49234;
    wire N__49233;
    wire N__49232;
    wire N__49231;
    wire N__49230;
    wire N__49229;
    wire N__49228;
    wire N__49227;
    wire N__49226;
    wire N__49225;
    wire N__49224;
    wire N__49223;
    wire N__49222;
    wire N__49221;
    wire N__49220;
    wire N__49219;
    wire N__49218;
    wire N__49217;
    wire N__49216;
    wire N__49215;
    wire N__49214;
    wire N__49213;
    wire N__49212;
    wire N__49211;
    wire N__49210;
    wire N__49209;
    wire N__49208;
    wire N__49207;
    wire N__49206;
    wire N__49205;
    wire N__49204;
    wire N__49203;
    wire N__49202;
    wire N__49201;
    wire N__49200;
    wire N__49199;
    wire N__49198;
    wire N__49197;
    wire N__49196;
    wire N__49195;
    wire N__49194;
    wire N__49193;
    wire N__49192;
    wire N__49191;
    wire N__49190;
    wire N__49189;
    wire N__49188;
    wire N__49187;
    wire N__49186;
    wire N__49185;
    wire N__49184;
    wire N__49183;
    wire N__49182;
    wire N__49181;
    wire N__49180;
    wire N__49179;
    wire N__49178;
    wire N__49177;
    wire N__49176;
    wire N__49175;
    wire N__49174;
    wire N__49173;
    wire N__49172;
    wire N__49171;
    wire N__49170;
    wire N__49169;
    wire N__49168;
    wire N__49167;
    wire N__49166;
    wire N__49165;
    wire N__49164;
    wire N__49163;
    wire N__49162;
    wire N__49161;
    wire N__49160;
    wire N__49159;
    wire N__49158;
    wire N__49157;
    wire N__49156;
    wire N__49155;
    wire N__49154;
    wire N__49153;
    wire N__49152;
    wire N__49151;
    wire N__49150;
    wire N__49149;
    wire N__49148;
    wire N__49147;
    wire N__49146;
    wire N__49145;
    wire N__49144;
    wire N__49143;
    wire N__49142;
    wire N__49141;
    wire N__49140;
    wire N__49139;
    wire N__49138;
    wire N__49137;
    wire N__49136;
    wire N__49135;
    wire N__49134;
    wire N__49133;
    wire N__49132;
    wire N__49131;
    wire N__49130;
    wire N__49129;
    wire N__49128;
    wire N__49127;
    wire N__49126;
    wire N__49125;
    wire N__49124;
    wire N__49123;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49119;
    wire N__49118;
    wire N__49117;
    wire N__49116;
    wire N__49115;
    wire N__49114;
    wire N__49113;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49108;
    wire N__49107;
    wire N__49106;
    wire N__49105;
    wire N__49104;
    wire N__49103;
    wire N__49102;
    wire N__49101;
    wire N__49100;
    wire N__49099;
    wire N__49098;
    wire N__49097;
    wire N__49096;
    wire N__49095;
    wire N__49094;
    wire N__49093;
    wire N__49092;
    wire N__49091;
    wire N__49090;
    wire N__49089;
    wire N__49088;
    wire N__48767;
    wire N__48764;
    wire N__48761;
    wire N__48760;
    wire N__48759;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48743;
    wire N__48740;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48732;
    wire N__48727;
    wire N__48724;
    wire N__48721;
    wire N__48716;
    wire N__48713;
    wire N__48712;
    wire N__48709;
    wire N__48708;
    wire N__48705;
    wire N__48702;
    wire N__48699;
    wire N__48694;
    wire N__48689;
    wire N__48686;
    wire N__48683;
    wire N__48682;
    wire N__48681;
    wire N__48678;
    wire N__48675;
    wire N__48672;
    wire N__48667;
    wire N__48662;
    wire N__48659;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48647;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48637;
    wire N__48632;
    wire N__48629;
    wire N__48628;
    wire N__48627;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48611;
    wire N__48608;
    wire N__48605;
    wire N__48604;
    wire N__48601;
    wire N__48598;
    wire N__48597;
    wire N__48592;
    wire N__48589;
    wire N__48586;
    wire N__48581;
    wire N__48578;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48567;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48551;
    wire N__48548;
    wire N__48545;
    wire N__48544;
    wire N__48541;
    wire N__48538;
    wire N__48537;
    wire N__48532;
    wire N__48529;
    wire N__48526;
    wire N__48521;
    wire N__48518;
    wire N__48517;
    wire N__48512;
    wire N__48511;
    wire N__48508;
    wire N__48505;
    wire N__48502;
    wire N__48497;
    wire N__48494;
    wire N__48493;
    wire N__48488;
    wire N__48487;
    wire N__48484;
    wire N__48481;
    wire N__48478;
    wire N__48473;
    wire N__48470;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48458;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48448;
    wire N__48443;
    wire N__48440;
    wire N__48439;
    wire N__48436;
    wire N__48433;
    wire N__48428;
    wire N__48427;
    wire N__48424;
    wire N__48421;
    wire N__48418;
    wire N__48413;
    wire N__48410;
    wire N__48409;
    wire N__48404;
    wire N__48403;
    wire N__48400;
    wire N__48397;
    wire N__48394;
    wire N__48389;
    wire N__48386;
    wire N__48383;
    wire N__48382;
    wire N__48379;
    wire N__48376;
    wire N__48375;
    wire N__48370;
    wire N__48367;
    wire N__48364;
    wire N__48359;
    wire N__48356;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48342;
    wire N__48337;
    wire N__48334;
    wire N__48331;
    wire N__48326;
    wire N__48323;
    wire N__48322;
    wire N__48319;
    wire N__48316;
    wire N__48315;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48299;
    wire N__48296;
    wire N__48293;
    wire N__48292;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48277;
    wire N__48276;
    wire N__48273;
    wire N__48270;
    wire N__48267;
    wire N__48264;
    wire N__48257;
    wire N__48254;
    wire N__48253;
    wire N__48252;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48236;
    wire N__48233;
    wire N__48232;
    wire N__48231;
    wire N__48226;
    wire N__48223;
    wire N__48220;
    wire N__48215;
    wire N__48212;
    wire N__48211;
    wire N__48208;
    wire N__48205;
    wire N__48202;
    wire N__48201;
    wire N__48196;
    wire N__48193;
    wire N__48190;
    wire N__48185;
    wire N__48182;
    wire N__48181;
    wire N__48178;
    wire N__48175;
    wire N__48172;
    wire N__48171;
    wire N__48166;
    wire N__48163;
    wire N__48160;
    wire N__48155;
    wire N__48152;
    wire N__48151;
    wire N__48148;
    wire N__48145;
    wire N__48140;
    wire N__48139;
    wire N__48136;
    wire N__48133;
    wire N__48130;
    wire N__48125;
    wire N__48122;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48110;
    wire N__48109;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48095;
    wire N__48092;
    wire N__48089;
    wire N__48088;
    wire N__48085;
    wire N__48082;
    wire N__48081;
    wire N__48076;
    wire N__48073;
    wire N__48070;
    wire N__48065;
    wire N__48062;
    wire N__48059;
    wire N__48056;
    wire N__48055;
    wire N__48052;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48042;
    wire N__48037;
    wire N__48034;
    wire N__48033;
    wire N__48030;
    wire N__48027;
    wire N__48024;
    wire N__48017;
    wire N__48014;
    wire N__48011;
    wire N__48010;
    wire N__48007;
    wire N__48004;
    wire N__48003;
    wire N__48000;
    wire N__47997;
    wire N__47994;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47984;
    wire N__47981;
    wire N__47972;
    wire N__47969;
    wire N__47968;
    wire N__47965;
    wire N__47962;
    wire N__47959;
    wire N__47956;
    wire N__47955;
    wire N__47952;
    wire N__47949;
    wire N__47946;
    wire N__47945;
    wire N__47942;
    wire N__47937;
    wire N__47934;
    wire N__47927;
    wire N__47924;
    wire N__47923;
    wire N__47920;
    wire N__47917;
    wire N__47914;
    wire N__47911;
    wire N__47910;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47879;
    wire N__47876;
    wire N__47875;
    wire N__47872;
    wire N__47869;
    wire N__47868;
    wire N__47863;
    wire N__47860;
    wire N__47859;
    wire N__47856;
    wire N__47853;
    wire N__47850;
    wire N__47843;
    wire N__47840;
    wire N__47837;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47827;
    wire N__47824;
    wire N__47823;
    wire N__47818;
    wire N__47815;
    wire N__47814;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47798;
    wire N__47795;
    wire N__47794;
    wire N__47793;
    wire N__47792;
    wire N__47791;
    wire N__47790;
    wire N__47789;
    wire N__47788;
    wire N__47771;
    wire N__47768;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47758;
    wire N__47757;
    wire N__47754;
    wire N__47751;
    wire N__47748;
    wire N__47745;
    wire N__47742;
    wire N__47739;
    wire N__47736;
    wire N__47731;
    wire N__47726;
    wire N__47723;
    wire N__47722;
    wire N__47719;
    wire N__47716;
    wire N__47713;
    wire N__47712;
    wire N__47709;
    wire N__47706;
    wire N__47703;
    wire N__47700;
    wire N__47693;
    wire N__47690;
    wire N__47689;
    wire N__47686;
    wire N__47685;
    wire N__47682;
    wire N__47679;
    wire N__47676;
    wire N__47675;
    wire N__47672;
    wire N__47667;
    wire N__47664;
    wire N__47661;
    wire N__47656;
    wire N__47651;
    wire N__47648;
    wire N__47645;
    wire N__47644;
    wire N__47643;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47615;
    wire N__47612;
    wire N__47603;
    wire N__47600;
    wire N__47599;
    wire N__47596;
    wire N__47595;
    wire N__47592;
    wire N__47589;
    wire N__47586;
    wire N__47581;
    wire N__47578;
    wire N__47577;
    wire N__47574;
    wire N__47571;
    wire N__47568;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47554;
    wire N__47551;
    wire N__47548;
    wire N__47545;
    wire N__47542;
    wire N__47541;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47519;
    wire N__47516;
    wire N__47513;
    wire N__47512;
    wire N__47509;
    wire N__47506;
    wire N__47503;
    wire N__47500;
    wire N__47495;
    wire N__47494;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47477;
    wire N__47474;
    wire N__47473;
    wire N__47470;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47460;
    wire N__47455;
    wire N__47452;
    wire N__47447;
    wire N__47446;
    wire N__47443;
    wire N__47440;
    wire N__47435;
    wire N__47432;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47421;
    wire N__47418;
    wire N__47415;
    wire N__47412;
    wire N__47409;
    wire N__47408;
    wire N__47405;
    wire N__47402;
    wire N__47399;
    wire N__47396;
    wire N__47387;
    wire N__47384;
    wire N__47383;
    wire N__47380;
    wire N__47377;
    wire N__47374;
    wire N__47371;
    wire N__47368;
    wire N__47367;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47355;
    wire N__47348;
    wire N__47345;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47328;
    wire N__47323;
    wire N__47322;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47306;
    wire N__47305;
    wire N__47302;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47284;
    wire N__47283;
    wire N__47278;
    wire N__47275;
    wire N__47272;
    wire N__47269;
    wire N__47264;
    wire N__47261;
    wire N__47260;
    wire N__47257;
    wire N__47256;
    wire N__47255;
    wire N__47252;
    wire N__47249;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47232;
    wire N__47227;
    wire N__47222;
    wire N__47219;
    wire N__47218;
    wire N__47217;
    wire N__47212;
    wire N__47209;
    wire N__47204;
    wire N__47201;
    wire N__47200;
    wire N__47197;
    wire N__47194;
    wire N__47189;
    wire N__47186;
    wire N__47183;
    wire N__47180;
    wire N__47179;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47169;
    wire N__47164;
    wire N__47163;
    wire N__47160;
    wire N__47157;
    wire N__47154;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47130;
    wire N__47129;
    wire N__47126;
    wire N__47123;
    wire N__47118;
    wire N__47113;
    wire N__47110;
    wire N__47105;
    wire N__47102;
    wire N__47099;
    wire N__47098;
    wire N__47095;
    wire N__47092;
    wire N__47091;
    wire N__47090;
    wire N__47085;
    wire N__47082;
    wire N__47079;
    wire N__47076;
    wire N__47073;
    wire N__47070;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47049;
    wire N__47048;
    wire N__47045;
    wire N__47042;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47028;
    wire N__47025;
    wire N__47020;
    wire N__47015;
    wire N__47012;
    wire N__47011;
    wire N__47008;
    wire N__47007;
    wire N__47004;
    wire N__47003;
    wire N__47000;
    wire N__46997;
    wire N__46994;
    wire N__46991;
    wire N__46988;
    wire N__46985;
    wire N__46980;
    wire N__46973;
    wire N__46970;
    wire N__46967;
    wire N__46964;
    wire N__46961;
    wire N__46958;
    wire N__46955;
    wire N__46952;
    wire N__46949;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46937;
    wire N__46934;
    wire N__46931;
    wire N__46930;
    wire N__46927;
    wire N__46924;
    wire N__46921;
    wire N__46918;
    wire N__46917;
    wire N__46914;
    wire N__46911;
    wire N__46908;
    wire N__46905;
    wire N__46904;
    wire N__46899;
    wire N__46896;
    wire N__46893;
    wire N__46890;
    wire N__46885;
    wire N__46880;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46868;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46856;
    wire N__46855;
    wire N__46852;
    wire N__46849;
    wire N__46844;
    wire N__46841;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46827;
    wire N__46822;
    wire N__46819;
    wire N__46818;
    wire N__46815;
    wire N__46812;
    wire N__46809;
    wire N__46806;
    wire N__46801;
    wire N__46796;
    wire N__46793;
    wire N__46790;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46782;
    wire N__46781;
    wire N__46778;
    wire N__46775;
    wire N__46772;
    wire N__46769;
    wire N__46766;
    wire N__46763;
    wire N__46760;
    wire N__46757;
    wire N__46754;
    wire N__46749;
    wire N__46746;
    wire N__46739;
    wire N__46736;
    wire N__46735;
    wire N__46732;
    wire N__46731;
    wire N__46728;
    wire N__46725;
    wire N__46722;
    wire N__46715;
    wire N__46714;
    wire N__46711;
    wire N__46708;
    wire N__46703;
    wire N__46700;
    wire N__46699;
    wire N__46696;
    wire N__46693;
    wire N__46690;
    wire N__46687;
    wire N__46686;
    wire N__46681;
    wire N__46678;
    wire N__46673;
    wire N__46670;
    wire N__46667;
    wire N__46664;
    wire N__46661;
    wire N__46660;
    wire N__46659;
    wire N__46658;
    wire N__46657;
    wire N__46654;
    wire N__46653;
    wire N__46652;
    wire N__46651;
    wire N__46650;
    wire N__46649;
    wire N__46648;
    wire N__46647;
    wire N__46646;
    wire N__46645;
    wire N__46644;
    wire N__46643;
    wire N__46642;
    wire N__46639;
    wire N__46638;
    wire N__46637;
    wire N__46636;
    wire N__46633;
    wire N__46632;
    wire N__46631;
    wire N__46630;
    wire N__46629;
    wire N__46628;
    wire N__46627;
    wire N__46626;
    wire N__46625;
    wire N__46624;
    wire N__46623;
    wire N__46622;
    wire N__46621;
    wire N__46614;
    wire N__46611;
    wire N__46610;
    wire N__46607;
    wire N__46606;
    wire N__46605;
    wire N__46604;
    wire N__46603;
    wire N__46602;
    wire N__46601;
    wire N__46600;
    wire N__46599;
    wire N__46598;
    wire N__46597;
    wire N__46596;
    wire N__46595;
    wire N__46594;
    wire N__46593;
    wire N__46592;
    wire N__46591;
    wire N__46590;
    wire N__46589;
    wire N__46588;
    wire N__46587;
    wire N__46584;
    wire N__46567;
    wire N__46566;
    wire N__46565;
    wire N__46564;
    wire N__46563;
    wire N__46562;
    wire N__46561;
    wire N__46560;
    wire N__46543;
    wire N__46528;
    wire N__46527;
    wire N__46526;
    wire N__46525;
    wire N__46524;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46513;
    wire N__46512;
    wire N__46511;
    wire N__46510;
    wire N__46509;
    wire N__46508;
    wire N__46507;
    wire N__46506;
    wire N__46505;
    wire N__46504;
    wire N__46501;
    wire N__46484;
    wire N__46481;
    wire N__46478;
    wire N__46477;
    wire N__46474;
    wire N__46473;
    wire N__46470;
    wire N__46469;
    wire N__46466;
    wire N__46463;
    wire N__46462;
    wire N__46459;
    wire N__46458;
    wire N__46455;
    wire N__46454;
    wire N__46451;
    wire N__46450;
    wire N__46449;
    wire N__46448;
    wire N__46447;
    wire N__46446;
    wire N__46445;
    wire N__46444;
    wire N__46443;
    wire N__46442;
    wire N__46441;
    wire N__46440;
    wire N__46439;
    wire N__46438;
    wire N__46435;
    wire N__46434;
    wire N__46431;
    wire N__46430;
    wire N__46427;
    wire N__46420;
    wire N__46417;
    wire N__46414;
    wire N__46399;
    wire N__46394;
    wire N__46389;
    wire N__46378;
    wire N__46377;
    wire N__46376;
    wire N__46375;
    wire N__46368;
    wire N__46367;
    wire N__46364;
    wire N__46363;
    wire N__46360;
    wire N__46359;
    wire N__46356;
    wire N__46355;
    wire N__46352;
    wire N__46349;
    wire N__46348;
    wire N__46345;
    wire N__46344;
    wire N__46341;
    wire N__46340;
    wire N__46337;
    wire N__46336;
    wire N__46333;
    wire N__46328;
    wire N__46313;
    wire N__46296;
    wire N__46293;
    wire N__46292;
    wire N__46289;
    wire N__46288;
    wire N__46285;
    wire N__46284;
    wire N__46281;
    wire N__46280;
    wire N__46277;
    wire N__46276;
    wire N__46273;
    wire N__46272;
    wire N__46269;
    wire N__46268;
    wire N__46265;
    wire N__46264;
    wire N__46261;
    wire N__46260;
    wire N__46257;
    wire N__46256;
    wire N__46253;
    wire N__46252;
    wire N__46239;
    wire N__46236;
    wire N__46229;
    wire N__46222;
    wire N__46215;
    wire N__46212;
    wire N__46195;
    wire N__46178;
    wire N__46169;
    wire N__46152;
    wire N__46135;
    wire N__46122;
    wire N__46119;
    wire N__46094;
    wire N__46093;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46058;
    wire N__46055;
    wire N__46052;
    wire N__46049;
    wire N__46046;
    wire N__46045;
    wire N__46042;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46032;
    wire N__46029;
    wire N__46026;
    wire N__46019;
    wire N__46016;
    wire N__46013;
    wire N__46010;
    wire N__46009;
    wire N__46008;
    wire N__46007;
    wire N__46006;
    wire N__46005;
    wire N__46004;
    wire N__46003;
    wire N__46002;
    wire N__46001;
    wire N__46000;
    wire N__45999;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45991;
    wire N__45988;
    wire N__45987;
    wire N__45986;
    wire N__45985;
    wire N__45984;
    wire N__45975;
    wire N__45966;
    wire N__45963;
    wire N__45962;
    wire N__45961;
    wire N__45960;
    wire N__45959;
    wire N__45958;
    wire N__45957;
    wire N__45956;
    wire N__45955;
    wire N__45952;
    wire N__45949;
    wire N__45944;
    wire N__45937;
    wire N__45926;
    wire N__45919;
    wire N__45918;
    wire N__45917;
    wire N__45916;
    wire N__45915;
    wire N__45914;
    wire N__45913;
    wire N__45912;
    wire N__45911;
    wire N__45910;
    wire N__45909;
    wire N__45908;
    wire N__45907;
    wire N__45900;
    wire N__45891;
    wire N__45888;
    wire N__45887;
    wire N__45886;
    wire N__45885;
    wire N__45884;
    wire N__45883;
    wire N__45882;
    wire N__45881;
    wire N__45880;
    wire N__45879;
    wire N__45878;
    wire N__45877;
    wire N__45876;
    wire N__45875;
    wire N__45874;
    wire N__45873;
    wire N__45872;
    wire N__45871;
    wire N__45870;
    wire N__45869;
    wire N__45856;
    wire N__45839;
    wire N__45838;
    wire N__45837;
    wire N__45836;
    wire N__45835;
    wire N__45834;
    wire N__45833;
    wire N__45832;
    wire N__45831;
    wire N__45830;
    wire N__45827;
    wire N__45826;
    wire N__45819;
    wire N__45814;
    wire N__45813;
    wire N__45810;
    wire N__45795;
    wire N__45780;
    wire N__45775;
    wire N__45768;
    wire N__45763;
    wire N__45752;
    wire N__45745;
    wire N__45738;
    wire N__45733;
    wire N__45730;
    wire N__45719;
    wire N__45716;
    wire N__45705;
    wire N__45702;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45685;
    wire N__45682;
    wire N__45679;
    wire N__45676;
    wire N__45673;
    wire N__45672;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45660;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45641;
    wire N__45638;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45615;
    wire N__45608;
    wire N__45605;
    wire N__45602;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45592;
    wire N__45591;
    wire N__45590;
    wire N__45589;
    wire N__45588;
    wire N__45587;
    wire N__45586;
    wire N__45585;
    wire N__45580;
    wire N__45573;
    wire N__45572;
    wire N__45569;
    wire N__45566;
    wire N__45561;
    wire N__45556;
    wire N__45553;
    wire N__45552;
    wire N__45551;
    wire N__45550;
    wire N__45549;
    wire N__45542;
    wire N__45537;
    wire N__45528;
    wire N__45527;
    wire N__45526;
    wire N__45525;
    wire N__45524;
    wire N__45523;
    wire N__45522;
    wire N__45521;
    wire N__45520;
    wire N__45519;
    wire N__45518;
    wire N__45517;
    wire N__45514;
    wire N__45509;
    wire N__45492;
    wire N__45489;
    wire N__45484;
    wire N__45473;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45456;
    wire N__45451;
    wire N__45446;
    wire N__45443;
    wire N__45440;
    wire N__45437;
    wire N__45434;
    wire N__45431;
    wire N__45428;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45416;
    wire N__45415;
    wire N__45412;
    wire N__45409;
    wire N__45408;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45374;
    wire N__45371;
    wire N__45368;
    wire N__45367;
    wire N__45366;
    wire N__45363;
    wire N__45360;
    wire N__45357;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45331;
    wire N__45328;
    wire N__45327;
    wire N__45322;
    wire N__45319;
    wire N__45316;
    wire N__45313;
    wire N__45310;
    wire N__45307;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45293;
    wire N__45290;
    wire N__45287;
    wire N__45286;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45276;
    wire N__45271;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45254;
    wire N__45251;
    wire N__45250;
    wire N__45249;
    wire N__45246;
    wire N__45243;
    wire N__45240;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45224;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45211;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45187;
    wire N__45184;
    wire N__45179;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45169;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45134;
    wire N__45131;
    wire N__45128;
    wire N__45127;
    wire N__45122;
    wire N__45119;
    wire N__45118;
    wire N__45117;
    wire N__45116;
    wire N__45115;
    wire N__45114;
    wire N__45113;
    wire N__45112;
    wire N__45111;
    wire N__45092;
    wire N__45089;
    wire N__45086;
    wire N__45085;
    wire N__45082;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45062;
    wire N__45059;
    wire N__45056;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45046;
    wire N__45043;
    wire N__45038;
    wire N__45035;
    wire N__45032;
    wire N__45029;
    wire N__45028;
    wire N__45025;
    wire N__45024;
    wire N__45023;
    wire N__45020;
    wire N__45017;
    wire N__45012;
    wire N__45009;
    wire N__45004;
    wire N__45003;
    wire N__44998;
    wire N__44995;
    wire N__44990;
    wire N__44989;
    wire N__44988;
    wire N__44987;
    wire N__44986;
    wire N__44985;
    wire N__44982;
    wire N__44981;
    wire N__44978;
    wire N__44977;
    wire N__44974;
    wire N__44973;
    wire N__44972;
    wire N__44971;
    wire N__44970;
    wire N__44969;
    wire N__44968;
    wire N__44967;
    wire N__44966;
    wire N__44965;
    wire N__44964;
    wire N__44963;
    wire N__44962;
    wire N__44961;
    wire N__44960;
    wire N__44959;
    wire N__44958;
    wire N__44953;
    wire N__44938;
    wire N__44937;
    wire N__44936;
    wire N__44935;
    wire N__44934;
    wire N__44931;
    wire N__44930;
    wire N__44927;
    wire N__44926;
    wire N__44923;
    wire N__44922;
    wire N__44919;
    wire N__44918;
    wire N__44917;
    wire N__44914;
    wire N__44913;
    wire N__44910;
    wire N__44909;
    wire N__44906;
    wire N__44905;
    wire N__44902;
    wire N__44895;
    wire N__44894;
    wire N__44893;
    wire N__44892;
    wire N__44891;
    wire N__44882;
    wire N__44877;
    wire N__44868;
    wire N__44851;
    wire N__44836;
    wire N__44835;
    wire N__44834;
    wire N__44833;
    wire N__44832;
    wire N__44831;
    wire N__44826;
    wire N__44817;
    wire N__44816;
    wire N__44815;
    wire N__44814;
    wire N__44813;
    wire N__44810;
    wire N__44801;
    wire N__44798;
    wire N__44793;
    wire N__44790;
    wire N__44787;
    wire N__44786;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44776;
    wire N__44771;
    wire N__44768;
    wire N__44763;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44747;
    wire N__44746;
    wire N__44735;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44721;
    wire N__44720;
    wire N__44717;
    wire N__44716;
    wire N__44715;
    wire N__44714;
    wire N__44713;
    wire N__44712;
    wire N__44711;
    wire N__44710;
    wire N__44709;
    wire N__44708;
    wire N__44705;
    wire N__44702;
    wire N__44695;
    wire N__44688;
    wire N__44685;
    wire N__44678;
    wire N__44669;
    wire N__44660;
    wire N__44651;
    wire N__44648;
    wire N__44645;
    wire N__44642;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44627;
    wire N__44624;
    wire N__44623;
    wire N__44620;
    wire N__44617;
    wire N__44612;
    wire N__44609;
    wire N__44606;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44598;
    wire N__44595;
    wire N__44592;
    wire N__44589;
    wire N__44586;
    wire N__44579;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44541;
    wire N__44538;
    wire N__44535;
    wire N__44532;
    wire N__44525;
    wire N__44522;
    wire N__44519;
    wire N__44516;
    wire N__44513;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44505;
    wire N__44500;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44480;
    wire N__44477;
    wire N__44474;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44466;
    wire N__44461;
    wire N__44458;
    wire N__44455;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44441;
    wire N__44438;
    wire N__44437;
    wire N__44436;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44420;
    wire N__44417;
    wire N__44416;
    wire N__44411;
    wire N__44410;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44396;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44386;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44364;
    wire N__44359;
    wire N__44356;
    wire N__44351;
    wire N__44348;
    wire N__44345;
    wire N__44342;
    wire N__44341;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44328;
    wire N__44321;
    wire N__44320;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44306;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44276;
    wire N__44273;
    wire N__44272;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44257;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44231;
    wire N__44228;
    wire N__44227;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44209;
    wire N__44204;
    wire N__44201;
    wire N__44200;
    wire N__44197;
    wire N__44192;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44177;
    wire N__44176;
    wire N__44173;
    wire N__44168;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44158;
    wire N__44153;
    wire N__44150;
    wire N__44147;
    wire N__44144;
    wire N__44141;
    wire N__44140;
    wire N__44139;
    wire N__44138;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44101;
    wire N__44098;
    wire N__44095;
    wire N__44090;
    wire N__44087;
    wire N__44086;
    wire N__44083;
    wire N__44080;
    wire N__44079;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44063;
    wire N__44060;
    wire N__44059;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44044;
    wire N__44041;
    wire N__44038;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44014;
    wire N__44011;
    wire N__44008;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43985;
    wire N__43984;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43969;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43951;
    wire N__43946;
    wire N__43943;
    wire N__43942;
    wire N__43939;
    wire N__43936;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43913;
    wire N__43912;
    wire N__43911;
    wire N__43906;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43880;
    wire N__43877;
    wire N__43876;
    wire N__43875;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43859;
    wire N__43856;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43841;
    wire N__43840;
    wire N__43839;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43827;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43811;
    wire N__43808;
    wire N__43805;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43790;
    wire N__43787;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43779;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43754;
    wire N__43751;
    wire N__43750;
    wire N__43749;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43723;
    wire N__43722;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43703;
    wire N__43702;
    wire N__43701;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43679;
    wire N__43676;
    wire N__43671;
    wire N__43668;
    wire N__43665;
    wire N__43662;
    wire N__43657;
    wire N__43652;
    wire N__43651;
    wire N__43650;
    wire N__43649;
    wire N__43646;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43624;
    wire N__43621;
    wire N__43618;
    wire N__43615;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43595;
    wire N__43592;
    wire N__43587;
    wire N__43580;
    wire N__43579;
    wire N__43574;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43559;
    wire N__43556;
    wire N__43555;
    wire N__43554;
    wire N__43551;
    wire N__43548;
    wire N__43545;
    wire N__43544;
    wire N__43541;
    wire N__43536;
    wire N__43533;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43500;
    wire N__43497;
    wire N__43490;
    wire N__43489;
    wire N__43488;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43476;
    wire N__43471;
    wire N__43468;
    wire N__43463;
    wire N__43460;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43449;
    wire N__43446;
    wire N__43443;
    wire N__43440;
    wire N__43437;
    wire N__43434;
    wire N__43427;
    wire N__43426;
    wire N__43425;
    wire N__43422;
    wire N__43417;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43391;
    wire N__43388;
    wire N__43387;
    wire N__43386;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43370;
    wire N__43369;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43351;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43334;
    wire N__43331;
    wire N__43330;
    wire N__43329;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43313;
    wire N__43310;
    wire N__43309;
    wire N__43308;
    wire N__43305;
    wire N__43300;
    wire N__43299;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43285;
    wire N__43280;
    wire N__43277;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43269;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43253;
    wire N__43252;
    wire N__43251;
    wire N__43248;
    wire N__43243;
    wire N__43240;
    wire N__43237;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43220;
    wire N__43217;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43205;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43190;
    wire N__43187;
    wire N__43184;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43176;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43150;
    wire N__43147;
    wire N__43146;
    wire N__43145;
    wire N__43142;
    wire N__43139;
    wire N__43134;
    wire N__43131;
    wire N__43124;
    wire N__43121;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43107;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43078;
    wire N__43077;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43065;
    wire N__43058;
    wire N__43055;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43047;
    wire N__43044;
    wire N__43041;
    wire N__43038;
    wire N__43033;
    wire N__43028;
    wire N__43025;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43017;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43005;
    wire N__42998;
    wire N__42995;
    wire N__42994;
    wire N__42993;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42977;
    wire N__42974;
    wire N__42973;
    wire N__42972;
    wire N__42971;
    wire N__42968;
    wire N__42963;
    wire N__42960;
    wire N__42953;
    wire N__42950;
    wire N__42949;
    wire N__42948;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42932;
    wire N__42929;
    wire N__42928;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42917;
    wire N__42914;
    wire N__42909;
    wire N__42906;
    wire N__42899;
    wire N__42896;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42888;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42872;
    wire N__42869;
    wire N__42868;
    wire N__42867;
    wire N__42864;
    wire N__42859;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42842;
    wire N__42839;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42827;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42812;
    wire N__42811;
    wire N__42808;
    wire N__42805;
    wire N__42804;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42788;
    wire N__42783;
    wire N__42780;
    wire N__42773;
    wire N__42770;
    wire N__42767;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42759;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42743;
    wire N__42742;
    wire N__42741;
    wire N__42738;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42726;
    wire N__42721;
    wire N__42718;
    wire N__42713;
    wire N__42710;
    wire N__42709;
    wire N__42706;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42691;
    wire N__42688;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42670;
    wire N__42667;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42649;
    wire N__42648;
    wire N__42643;
    wire N__42640;
    wire N__42635;
    wire N__42632;
    wire N__42631;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42613;
    wire N__42612;
    wire N__42607;
    wire N__42604;
    wire N__42599;
    wire N__42596;
    wire N__42595;
    wire N__42594;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42578;
    wire N__42575;
    wire N__42574;
    wire N__42573;
    wire N__42570;
    wire N__42565;
    wire N__42560;
    wire N__42557;
    wire N__42556;
    wire N__42553;
    wire N__42550;
    wire N__42545;
    wire N__42542;
    wire N__42541;
    wire N__42540;
    wire N__42535;
    wire N__42532;
    wire N__42529;
    wire N__42524;
    wire N__42521;
    wire N__42520;
    wire N__42517;
    wire N__42514;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42503;
    wire N__42500;
    wire N__42497;
    wire N__42494;
    wire N__42491;
    wire N__42482;
    wire N__42479;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42471;
    wire N__42466;
    wire N__42463;
    wire N__42460;
    wire N__42455;
    wire N__42454;
    wire N__42451;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42433;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42416;
    wire N__42413;
    wire N__42412;
    wire N__42409;
    wire N__42406;
    wire N__42405;
    wire N__42400;
    wire N__42397;
    wire N__42394;
    wire N__42389;
    wire N__42388;
    wire N__42385;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42369;
    wire N__42364;
    wire N__42363;
    wire N__42358;
    wire N__42355;
    wire N__42350;
    wire N__42347;
    wire N__42346;
    wire N__42341;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42326;
    wire N__42323;
    wire N__42322;
    wire N__42319;
    wire N__42318;
    wire N__42317;
    wire N__42314;
    wire N__42311;
    wire N__42308;
    wire N__42305;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42289;
    wire N__42286;
    wire N__42283;
    wire N__42282;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42266;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42254;
    wire N__42251;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42224;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42197;
    wire N__42194;
    wire N__42191;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42179;
    wire N__42178;
    wire N__42177;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42113;
    wire N__42110;
    wire N__42107;
    wire N__42104;
    wire N__42101;
    wire N__42098;
    wire N__42095;
    wire N__42092;
    wire N__42089;
    wire N__42086;
    wire N__42083;
    wire N__42080;
    wire N__42079;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42062;
    wire N__42059;
    wire N__42056;
    wire N__42053;
    wire N__42052;
    wire N__42051;
    wire N__42048;
    wire N__42045;
    wire N__42042;
    wire N__42035;
    wire N__42032;
    wire N__42029;
    wire N__42026;
    wire N__42023;
    wire N__42022;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__41999;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41983;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41963;
    wire N__41960;
    wire N__41957;
    wire N__41954;
    wire N__41951;
    wire N__41948;
    wire N__41947;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41918;
    wire N__41917;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41885;
    wire N__41882;
    wire N__41879;
    wire N__41876;
    wire N__41873;
    wire N__41872;
    wire N__41871;
    wire N__41870;
    wire N__41869;
    wire N__41868;
    wire N__41867;
    wire N__41866;
    wire N__41865;
    wire N__41864;
    wire N__41863;
    wire N__41862;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41838;
    wire N__41837;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41827;
    wire N__41826;
    wire N__41825;
    wire N__41824;
    wire N__41823;
    wire N__41822;
    wire N__41815;
    wire N__41812;
    wire N__41811;
    wire N__41810;
    wire N__41809;
    wire N__41808;
    wire N__41807;
    wire N__41806;
    wire N__41805;
    wire N__41804;
    wire N__41803;
    wire N__41802;
    wire N__41801;
    wire N__41800;
    wire N__41797;
    wire N__41792;
    wire N__41789;
    wire N__41778;
    wire N__41773;
    wire N__41756;
    wire N__41747;
    wire N__41744;
    wire N__41737;
    wire N__41734;
    wire N__41729;
    wire N__41720;
    wire N__41717;
    wire N__41716;
    wire N__41715;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41699;
    wire N__41696;
    wire N__41693;
    wire N__41690;
    wire N__41687;
    wire N__41684;
    wire N__41681;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41669;
    wire N__41666;
    wire N__41663;
    wire N__41660;
    wire N__41657;
    wire N__41654;
    wire N__41651;
    wire N__41648;
    wire N__41645;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41615;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41600;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41563;
    wire N__41562;
    wire N__41561;
    wire N__41560;
    wire N__41559;
    wire N__41558;
    wire N__41557;
    wire N__41556;
    wire N__41555;
    wire N__41554;
    wire N__41553;
    wire N__41552;
    wire N__41551;
    wire N__41550;
    wire N__41549;
    wire N__41548;
    wire N__41547;
    wire N__41546;
    wire N__41545;
    wire N__41544;
    wire N__41543;
    wire N__41542;
    wire N__41541;
    wire N__41540;
    wire N__41539;
    wire N__41538;
    wire N__41537;
    wire N__41536;
    wire N__41535;
    wire N__41526;
    wire N__41517;
    wire N__41508;
    wire N__41499;
    wire N__41490;
    wire N__41481;
    wire N__41476;
    wire N__41467;
    wire N__41462;
    wire N__41459;
    wire N__41448;
    wire N__41441;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41431;
    wire N__41430;
    wire N__41427;
    wire N__41424;
    wire N__41421;
    wire N__41420;
    wire N__41417;
    wire N__41414;
    wire N__41411;
    wire N__41408;
    wire N__41405;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41385;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41331;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41300;
    wire N__41297;
    wire N__41294;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41273;
    wire N__41270;
    wire N__41267;
    wire N__41264;
    wire N__41261;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41246;
    wire N__41243;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41222;
    wire N__41219;
    wire N__41216;
    wire N__41213;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41170;
    wire N__41167;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41090;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41059;
    wire N__41056;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41039;
    wire N__41036;
    wire N__41033;
    wire N__41030;
    wire N__41027;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__41001;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40972;
    wire N__40969;
    wire N__40966;
    wire N__40961;
    wire N__40960;
    wire N__40957;
    wire N__40954;
    wire N__40953;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40937;
    wire N__40936;
    wire N__40933;
    wire N__40928;
    wire N__40927;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40913;
    wire N__40910;
    wire N__40907;
    wire N__40904;
    wire N__40901;
    wire N__40898;
    wire N__40895;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40883;
    wire N__40880;
    wire N__40877;
    wire N__40876;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40864;
    wire N__40861;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40844;
    wire N__40843;
    wire N__40840;
    wire N__40837;
    wire N__40836;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40805;
    wire N__40802;
    wire N__40799;
    wire N__40796;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40757;
    wire N__40754;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40742;
    wire N__40739;
    wire N__40736;
    wire N__40733;
    wire N__40732;
    wire N__40729;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40712;
    wire N__40709;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40695;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40679;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40667;
    wire N__40666;
    wire N__40663;
    wire N__40662;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40643;
    wire N__40640;
    wire N__40637;
    wire N__40634;
    wire N__40631;
    wire N__40628;
    wire N__40627;
    wire N__40626;
    wire N__40619;
    wire N__40616;
    wire N__40613;
    wire N__40610;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40586;
    wire N__40583;
    wire N__40582;
    wire N__40577;
    wire N__40574;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40550;
    wire N__40547;
    wire N__40544;
    wire N__40541;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40529;
    wire N__40526;
    wire N__40523;
    wire N__40520;
    wire N__40517;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40489;
    wire N__40488;
    wire N__40483;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40473;
    wire N__40470;
    wire N__40467;
    wire N__40464;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40450;
    wire N__40447;
    wire N__40446;
    wire N__40445;
    wire N__40440;
    wire N__40435;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40417;
    wire N__40414;
    wire N__40411;
    wire N__40406;
    wire N__40405;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40364;
    wire N__40361;
    wire N__40358;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40334;
    wire N__40333;
    wire N__40328;
    wire N__40327;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40313;
    wire N__40310;
    wire N__40309;
    wire N__40304;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40289;
    wire N__40286;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40265;
    wire N__40264;
    wire N__40259;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40249;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40234;
    wire N__40229;
    wire N__40226;
    wire N__40225;
    wire N__40220;
    wire N__40217;
    wire N__40216;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40168;
    wire N__40165;
    wire N__40164;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40148;
    wire N__40147;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40135;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40118;
    wire N__40115;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40103;
    wire N__40102;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40085;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40070;
    wire N__40069;
    wire N__40064;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40049;
    wire N__40046;
    wire N__40045;
    wire N__40040;
    wire N__40037;
    wire N__40036;
    wire N__40033;
    wire N__40028;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40013;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__40000;
    wire N__39997;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39980;
    wire N__39979;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39956;
    wire N__39953;
    wire N__39950;
    wire N__39947;
    wire N__39944;
    wire N__39943;
    wire N__39938;
    wire N__39937;
    wire N__39934;
    wire N__39931;
    wire N__39928;
    wire N__39923;
    wire N__39920;
    wire N__39919;
    wire N__39914;
    wire N__39913;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39899;
    wire N__39898;
    wire N__39893;
    wire N__39890;
    wire N__39887;
    wire N__39884;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39874;
    wire N__39871;
    wire N__39868;
    wire N__39863;
    wire N__39860;
    wire N__39859;
    wire N__39854;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39844;
    wire N__39839;
    wire N__39836;
    wire N__39835;
    wire N__39834;
    wire N__39831;
    wire N__39826;
    wire N__39821;
    wire N__39820;
    wire N__39819;
    wire N__39816;
    wire N__39811;
    wire N__39806;
    wire N__39803;
    wire N__39800;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39772;
    wire N__39767;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39757;
    wire N__39752;
    wire N__39751;
    wire N__39748;
    wire N__39743;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39728;
    wire N__39725;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39712;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39700;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39688;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39667;
    wire N__39666;
    wire N__39663;
    wire N__39658;
    wire N__39653;
    wire N__39652;
    wire N__39649;
    wire N__39648;
    wire N__39645;
    wire N__39640;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39610;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39598;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39581;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39571;
    wire N__39568;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39551;
    wire N__39550;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39542;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39518;
    wire N__39515;
    wire N__39506;
    wire N__39505;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39451;
    wire N__39450;
    wire N__39447;
    wire N__39442;
    wire N__39439;
    wire N__39438;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39426;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39397;
    wire N__39396;
    wire N__39391;
    wire N__39388;
    wire N__39385;
    wire N__39380;
    wire N__39377;
    wire N__39376;
    wire N__39371;
    wire N__39370;
    wire N__39367;
    wire N__39364;
    wire N__39361;
    wire N__39356;
    wire N__39353;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39341;
    wire N__39340;
    wire N__39335;
    wire N__39332;
    wire N__39329;
    wire N__39326;
    wire N__39323;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39293;
    wire N__39292;
    wire N__39289;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39272;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39257;
    wire N__39256;
    wire N__39255;
    wire N__39252;
    wire N__39251;
    wire N__39246;
    wire N__39241;
    wire N__39238;
    wire N__39233;
    wire N__39232;
    wire N__39229;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39214;
    wire N__39211;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39194;
    wire N__39191;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39125;
    wire N__39122;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39080;
    wire N__39077;
    wire N__39074;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39062;
    wire N__39059;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38969;
    wire N__38966;
    wire N__38963;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38939;
    wire N__38936;
    wire N__38933;
    wire N__38930;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38819;
    wire N__38816;
    wire N__38813;
    wire N__38810;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38798;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38735;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38699;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38663;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38648;
    wire N__38645;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38555;
    wire N__38552;
    wire N__38549;
    wire N__38546;
    wire N__38543;
    wire N__38540;
    wire N__38537;
    wire N__38534;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38420;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38399;
    wire N__38396;
    wire N__38393;
    wire N__38392;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38333;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38312;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38270;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38249;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38228;
    wire N__38225;
    wire N__38222;
    wire N__38219;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38189;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38177;
    wire N__38174;
    wire N__38171;
    wire N__38168;
    wire N__38165;
    wire N__38162;
    wire N__38161;
    wire N__38158;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38142;
    wire N__38137;
    wire N__38132;
    wire N__38129;
    wire N__38126;
    wire N__38123;
    wire N__38120;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38108;
    wire N__38105;
    wire N__38102;
    wire N__38099;
    wire N__38096;
    wire N__38093;
    wire N__38090;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38075;
    wire N__38072;
    wire N__38069;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38000;
    wire N__37997;
    wire N__37994;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37955;
    wire N__37952;
    wire N__37949;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37937;
    wire N__37936;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37918;
    wire N__37913;
    wire N__37912;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37889;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37877;
    wire N__37876;
    wire N__37873;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37856;
    wire N__37855;
    wire N__37852;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37822;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37802;
    wire N__37799;
    wire N__37798;
    wire N__37795;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37772;
    wire N__37769;
    wire N__37768;
    wire N__37765;
    wire N__37764;
    wire N__37761;
    wire N__37756;
    wire N__37751;
    wire N__37748;
    wire N__37747;
    wire N__37746;
    wire N__37743;
    wire N__37738;
    wire N__37733;
    wire N__37730;
    wire N__37727;
    wire N__37724;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37712;
    wire N__37709;
    wire N__37708;
    wire N__37705;
    wire N__37702;
    wire N__37697;
    wire N__37694;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37682;
    wire N__37679;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37657;
    wire N__37654;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37637;
    wire N__37634;
    wire N__37633;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37616;
    wire N__37613;
    wire N__37612;
    wire N__37609;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37586;
    wire N__37583;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37571;
    wire N__37568;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37556;
    wire N__37553;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37541;
    wire N__37538;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37526;
    wire N__37523;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37511;
    wire N__37508;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37496;
    wire N__37493;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37481;
    wire N__37478;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37466;
    wire N__37463;
    wire N__37462;
    wire N__37461;
    wire N__37460;
    wire N__37457;
    wire N__37452;
    wire N__37449;
    wire N__37442;
    wire N__37441;
    wire N__37440;
    wire N__37439;
    wire N__37436;
    wire N__37431;
    wire N__37428;
    wire N__37421;
    wire N__37420;
    wire N__37417;
    wire N__37416;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37363;
    wire N__37360;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37345;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37319;
    wire N__37318;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37304;
    wire N__37301;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36920;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36880;
    wire N__36879;
    wire N__36878;
    wire N__36877;
    wire N__36876;
    wire N__36875;
    wire N__36874;
    wire N__36871;
    wire N__36870;
    wire N__36869;
    wire N__36868;
    wire N__36867;
    wire N__36866;
    wire N__36865;
    wire N__36864;
    wire N__36863;
    wire N__36862;
    wire N__36861;
    wire N__36860;
    wire N__36859;
    wire N__36858;
    wire N__36857;
    wire N__36856;
    wire N__36855;
    wire N__36854;
    wire N__36853;
    wire N__36852;
    wire N__36851;
    wire N__36844;
    wire N__36835;
    wire N__36834;
    wire N__36833;
    wire N__36832;
    wire N__36831;
    wire N__36828;
    wire N__36819;
    wire N__36810;
    wire N__36801;
    wire N__36792;
    wire N__36783;
    wire N__36778;
    wire N__36769;
    wire N__36766;
    wire N__36761;
    wire N__36750;
    wire N__36747;
    wire N__36742;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36728;
    wire N__36725;
    wire N__36724;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36701;
    wire N__36700;
    wire N__36697;
    wire N__36696;
    wire N__36693;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36682;
    wire N__36679;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36655;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36637;
    wire N__36632;
    wire N__36631;
    wire N__36628;
    wire N__36625;
    wire N__36622;
    wire N__36617;
    wire N__36614;
    wire N__36613;
    wire N__36612;
    wire N__36607;
    wire N__36604;
    wire N__36601;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36487;
    wire N__36484;
    wire N__36481;
    wire N__36478;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36460;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36443;
    wire N__36442;
    wire N__36437;
    wire N__36434;
    wire N__36433;
    wire N__36430;
    wire N__36427;
    wire N__36422;
    wire N__36419;
    wire N__36418;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36397;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36371;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36343;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36320;
    wire N__36317;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36200;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36157;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36147;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36113;
    wire N__36110;
    wire N__36109;
    wire N__36108;
    wire N__36105;
    wire N__36100;
    wire N__36097;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35995;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35966;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35958;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35915;
    wire N__35912;
    wire N__35911;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35894;
    wire N__35891;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35887;
    wire N__35886;
    wire N__35883;
    wire N__35878;
    wire N__35875;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35825;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35805;
    wire N__35802;
    wire N__35799;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35704;
    wire N__35701;
    wire N__35700;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35687;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35671;
    wire N__35668;
    wire N__35667;
    wire N__35664;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35646;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35628;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35546;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35531;
    wire N__35528;
    wire N__35527;
    wire N__35526;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35488;
    wire N__35483;
    wire N__35480;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35463;
    wire N__35460;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35441;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35430;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35418;
    wire N__35415;
    wire N__35410;
    wire N__35407;
    wire N__35402;
    wire N__35399;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35391;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35375;
    wire N__35374;
    wire N__35371;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35303;
    wire N__35300;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35292;
    wire N__35287;
    wire N__35284;
    wire N__35281;
    wire N__35276;
    wire N__35275;
    wire N__35272;
    wire N__35271;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35259;
    wire N__35256;
    wire N__35251;
    wire N__35248;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35219;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35207;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35192;
    wire N__35191;
    wire N__35190;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35180;
    wire N__35177;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35149;
    wire N__35148;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35135;
    wire N__35132;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35105;
    wire N__35104;
    wire N__35101;
    wire N__35100;
    wire N__35099;
    wire N__35096;
    wire N__35093;
    wire N__35090;
    wire N__35087;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35056;
    wire N__35053;
    wire N__35048;
    wire N__35043;
    wire N__35036;
    wire N__35035;
    wire N__35030;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35015;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35007;
    wire N__35002;
    wire N__34999;
    wire N__34998;
    wire N__34993;
    wire N__34990;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34943;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34935;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34900;
    wire N__34895;
    wire N__34892;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34863;
    wire N__34856;
    wire N__34853;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34845;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34830;
    wire N__34825;
    wire N__34822;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34800;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34784;
    wire N__34781;
    wire N__34778;
    wire N__34777;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34766;
    wire N__34759;
    wire N__34756;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34734;
    wire N__34729;
    wire N__34726;
    wire N__34723;
    wire N__34718;
    wire N__34717;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34706;
    wire N__34703;
    wire N__34698;
    wire N__34695;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34662;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34646;
    wire N__34645;
    wire N__34644;
    wire N__34641;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34617;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34601;
    wire N__34598;
    wire N__34597;
    wire N__34592;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34577;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34562;
    wire N__34559;
    wire N__34556;
    wire N__34553;
    wire N__34546;
    wire N__34543;
    wire N__34538;
    wire N__34535;
    wire N__34534;
    wire N__34529;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34509;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34472;
    wire N__34469;
    wire N__34468;
    wire N__34467;
    wire N__34464;
    wire N__34459;
    wire N__34458;
    wire N__34453;
    wire N__34450;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34408;
    wire N__34405;
    wire N__34400;
    wire N__34397;
    wire N__34396;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34385;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34348;
    wire N__34347;
    wire N__34344;
    wire N__34341;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34327;
    wire N__34324;
    wire N__34319;
    wire N__34316;
    wire N__34315;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34260;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34244;
    wire N__34243;
    wire N__34240;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34230;
    wire N__34229;
    wire N__34226;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34210;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34191;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34175;
    wire N__34174;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34144;
    wire N__34141;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34122;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34106;
    wire N__34103;
    wire N__34102;
    wire N__34101;
    wire N__34100;
    wire N__34097;
    wire N__34092;
    wire N__34089;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34062;
    wire N__34057;
    wire N__34054;
    wire N__34051;
    wire N__34046;
    wire N__34045;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34030;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33990;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33974;
    wire N__33971;
    wire N__33970;
    wire N__33969;
    wire N__33966;
    wire N__33961;
    wire N__33960;
    wire N__33955;
    wire N__33952;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33908;
    wire N__33907;
    wire N__33904;
    wire N__33903;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33874;
    wire N__33869;
    wire N__33866;
    wire N__33865;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33844;
    wire N__33839;
    wire N__33838;
    wire N__33835;
    wire N__33834;
    wire N__33831;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33794;
    wire N__33791;
    wire N__33790;
    wire N__33785;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33770;
    wire N__33769;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33729;
    wire N__33724;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33705;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33689;
    wire N__33688;
    wire N__33687;
    wire N__33684;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33652;
    wire N__33647;
    wire N__33644;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33633;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33617;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33609;
    wire N__33608;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33580;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33561;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33545;
    wire N__33544;
    wire N__33539;
    wire N__33538;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33511;
    wire N__33506;
    wire N__33503;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33491;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33476;
    wire N__33475;
    wire N__33474;
    wire N__33471;
    wire N__33466;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33417;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33385;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33353;
    wire N__33352;
    wire N__33351;
    wire N__33348;
    wire N__33345;
    wire N__33342;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33211;
    wire N__33208;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33056;
    wire N__33053;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33041;
    wire N__33038;
    wire N__33035;
    wire N__33032;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32935;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32840;
    wire N__32837;
    wire N__32834;
    wire N__32831;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32791;
    wire N__32790;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32774;
    wire N__32771;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32746;
    wire N__32741;
    wire N__32738;
    wire N__32737;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32726;
    wire N__32725;
    wire N__32724;
    wire N__32723;
    wire N__32722;
    wire N__32721;
    wire N__32716;
    wire N__32715;
    wire N__32714;
    wire N__32713;
    wire N__32712;
    wire N__32711;
    wire N__32710;
    wire N__32709;
    wire N__32708;
    wire N__32707;
    wire N__32706;
    wire N__32705;
    wire N__32704;
    wire N__32703;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32692;
    wire N__32691;
    wire N__32690;
    wire N__32689;
    wire N__32688;
    wire N__32687;
    wire N__32680;
    wire N__32679;
    wire N__32676;
    wire N__32675;
    wire N__32674;
    wire N__32673;
    wire N__32672;
    wire N__32671;
    wire N__32670;
    wire N__32669;
    wire N__32668;
    wire N__32667;
    wire N__32666;
    wire N__32665;
    wire N__32662;
    wire N__32653;
    wire N__32644;
    wire N__32635;
    wire N__32632;
    wire N__32631;
    wire N__32628;
    wire N__32627;
    wire N__32620;
    wire N__32611;
    wire N__32608;
    wire N__32605;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32587;
    wire N__32580;
    wire N__32571;
    wire N__32564;
    wire N__32561;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32534;
    wire N__32529;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32507;
    wire N__32500;
    wire N__32495;
    wire N__32490;
    wire N__32477;
    wire N__32474;
    wire N__32473;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32458;
    wire N__32453;
    wire N__32450;
    wire N__32449;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32426;
    wire N__32425;
    wire N__32424;
    wire N__32423;
    wire N__32422;
    wire N__32421;
    wire N__32420;
    wire N__32419;
    wire N__32418;
    wire N__32417;
    wire N__32416;
    wire N__32415;
    wire N__32414;
    wire N__32413;
    wire N__32412;
    wire N__32411;
    wire N__32410;
    wire N__32409;
    wire N__32408;
    wire N__32407;
    wire N__32406;
    wire N__32405;
    wire N__32404;
    wire N__32403;
    wire N__32402;
    wire N__32401;
    wire N__32400;
    wire N__32399;
    wire N__32398;
    wire N__32397;
    wire N__32396;
    wire N__32395;
    wire N__32394;
    wire N__32393;
    wire N__32392;
    wire N__32387;
    wire N__32380;
    wire N__32373;
    wire N__32368;
    wire N__32363;
    wire N__32362;
    wire N__32361;
    wire N__32360;
    wire N__32359;
    wire N__32358;
    wire N__32357;
    wire N__32356;
    wire N__32355;
    wire N__32354;
    wire N__32353;
    wire N__32352;
    wire N__32351;
    wire N__32350;
    wire N__32349;
    wire N__32348;
    wire N__32347;
    wire N__32346;
    wire N__32345;
    wire N__32344;
    wire N__32341;
    wire N__32340;
    wire N__32339;
    wire N__32338;
    wire N__32337;
    wire N__32336;
    wire N__32335;
    wire N__32334;
    wire N__32333;
    wire N__32332;
    wire N__32331;
    wire N__32330;
    wire N__32329;
    wire N__32328;
    wire N__32327;
    wire N__32326;
    wire N__32325;
    wire N__32324;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32309;
    wire N__32308;
    wire N__32307;
    wire N__32306;
    wire N__32305;
    wire N__32304;
    wire N__32303;
    wire N__32300;
    wire N__32291;
    wire N__32278;
    wire N__32269;
    wire N__32264;
    wire N__32253;
    wire N__32242;
    wire N__32239;
    wire N__32228;
    wire N__32217;
    wire N__32210;
    wire N__32207;
    wire N__32200;
    wire N__32191;
    wire N__32190;
    wire N__32189;
    wire N__32188;
    wire N__32187;
    wire N__32186;
    wire N__32185;
    wire N__32184;
    wire N__32171;
    wire N__32170;
    wire N__32169;
    wire N__32168;
    wire N__32167;
    wire N__32166;
    wire N__32165;
    wire N__32164;
    wire N__32161;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32143;
    wire N__32128;
    wire N__32115;
    wire N__32112;
    wire N__32107;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32079;
    wire N__32076;
    wire N__32067;
    wire N__32062;
    wire N__32059;
    wire N__32054;
    wire N__32051;
    wire N__32048;
    wire N__32041;
    wire N__32038;
    wire N__32033;
    wire N__32006;
    wire N__32003;
    wire N__32002;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31979;
    wire N__31976;
    wire N__31975;
    wire N__31972;
    wire N__31969;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31954;
    wire N__31951;
    wire N__31950;
    wire N__31947;
    wire N__31946;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31925;
    wire N__31922;
    wire N__31913;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31901;
    wire N__31900;
    wire N__31897;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31874;
    wire N__31871;
    wire N__31870;
    wire N__31867;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31852;
    wire N__31847;
    wire N__31844;
    wire N__31843;
    wire N__31838;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31823;
    wire N__31820;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31806;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31790;
    wire N__31787;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31779;
    wire N__31774;
    wire N__31771;
    wire N__31768;
    wire N__31763;
    wire N__31760;
    wire N__31759;
    wire N__31754;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31739;
    wire N__31736;
    wire N__31733;
    wire N__31732;
    wire N__31731;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31715;
    wire N__31712;
    wire N__31711;
    wire N__31710;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31694;
    wire N__31691;
    wire N__31688;
    wire N__31687;
    wire N__31686;
    wire N__31681;
    wire N__31678;
    wire N__31675;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31579;
    wire N__31574;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31559;
    wire N__31556;
    wire N__31555;
    wire N__31554;
    wire N__31549;
    wire N__31546;
    wire N__31543;
    wire N__31538;
    wire N__31535;
    wire N__31534;
    wire N__31529;
    wire N__31526;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31511;
    wire N__31508;
    wire N__31507;
    wire N__31504;
    wire N__31499;
    wire N__31496;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31313;
    wire N__31310;
    wire N__31309;
    wire N__31306;
    wire N__31305;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31289;
    wire N__31286;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31235;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31218;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31171;
    wire N__31168;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31072;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31049;
    wire N__31048;
    wire N__31047;
    wire N__31046;
    wire N__31043;
    wire N__31036;
    wire N__31033;
    wire N__31028;
    wire N__31027;
    wire N__31024;
    wire N__31023;
    wire N__31022;
    wire N__31015;
    wire N__31012;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30988;
    wire N__30985;
    wire N__30982;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30952;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30851;
    wire N__30848;
    wire N__30845;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30545;
    wire N__30542;
    wire N__30539;
    wire N__30536;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30425;
    wire N__30422;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30401;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30302;
    wire N__30299;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30286;
    wire N__30283;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30236;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30200;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30074;
    wire N__30071;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30037;
    wire N__30034;
    wire N__30033;
    wire N__30028;
    wire N__30025;
    wire N__30020;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30008;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29996;
    wire N__29995;
    wire N__29994;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29935;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29925;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29902;
    wire N__29899;
    wire N__29896;
    wire N__29891;
    wire N__29888;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29880;
    wire N__29875;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29858;
    wire N__29857;
    wire N__29856;
    wire N__29853;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29813;
    wire N__29812;
    wire N__29809;
    wire N__29808;
    wire N__29807;
    wire N__29804;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29786;
    wire N__29785;
    wire N__29784;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29772;
    wire N__29765;
    wire N__29764;
    wire N__29763;
    wire N__29762;
    wire N__29753;
    wire N__29752;
    wire N__29751;
    wire N__29750;
    wire N__29749;
    wire N__29748;
    wire N__29747;
    wire N__29746;
    wire N__29745;
    wire N__29744;
    wire N__29743;
    wire N__29742;
    wire N__29741;
    wire N__29740;
    wire N__29739;
    wire N__29738;
    wire N__29737;
    wire N__29736;
    wire N__29735;
    wire N__29734;
    wire N__29733;
    wire N__29732;
    wire N__29731;
    wire N__29728;
    wire N__29719;
    wire N__29710;
    wire N__29709;
    wire N__29708;
    wire N__29707;
    wire N__29706;
    wire N__29701;
    wire N__29692;
    wire N__29683;
    wire N__29674;
    wire N__29667;
    wire N__29658;
    wire N__29645;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29633;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29577;
    wire N__29572;
    wire N__29571;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29559;
    wire N__29552;
    wire N__29549;
    wire N__29548;
    wire N__29545;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29470;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29455;
    wire N__29454;
    wire N__29453;
    wire N__29450;
    wire N__29443;
    wire N__29438;
    wire N__29435;
    wire N__29432;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29416;
    wire N__29413;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29356;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29344;
    wire N__29341;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29324;
    wire N__29323;
    wire N__29318;
    wire N__29315;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29293;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29272;
    wire N__29271;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29259;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29240;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29229;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29204;
    wire N__29201;
    wire N__29200;
    wire N__29197;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29180;
    wire N__29179;
    wire N__29176;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29119;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29105;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29087;
    wire N__29086;
    wire N__29085;
    wire N__29080;
    wire N__29077;
    wire N__29072;
    wire N__29069;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29024;
    wire N__29021;
    wire N__29020;
    wire N__29019;
    wire N__29016;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29003;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28975;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28958;
    wire N__28957;
    wire N__28954;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28937;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28922;
    wire N__28921;
    wire N__28920;
    wire N__28919;
    wire N__28918;
    wire N__28917;
    wire N__28916;
    wire N__28915;
    wire N__28914;
    wire N__28913;
    wire N__28912;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28882;
    wire N__28881;
    wire N__28878;
    wire N__28873;
    wire N__28868;
    wire N__28867;
    wire N__28866;
    wire N__28863;
    wire N__28862;
    wire N__28857;
    wire N__28852;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28795;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28767;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28755;
    wire N__28748;
    wire N__28747;
    wire N__28744;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28720;
    wire N__28717;
    wire N__28712;
    wire N__28711;
    wire N__28706;
    wire N__28703;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28667;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28655;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28643;
    wire N__28640;
    wire N__28639;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28582;
    wire N__28579;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28562;
    wire N__28561;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28544;
    wire N__28543;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28528;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28507;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28421;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28402;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28370;
    wire N__28369;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28045;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28028;
    wire N__28027;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28010;
    wire N__28009;
    wire N__28004;
    wire N__28001;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27989;
    wire N__27988;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27910;
    wire N__27905;
    wire N__27902;
    wire N__27901;
    wire N__27898;
    wire N__27893;
    wire N__27890;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27860;
    wire N__27859;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27844;
    wire N__27839;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27802;
    wire N__27797;
    wire N__27794;
    wire N__27793;
    wire N__27788;
    wire N__27785;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27763;
    wire N__27758;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27698;
    wire N__27695;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27683;
    wire N__27680;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27668;
    wire N__27665;
    wire N__27664;
    wire N__27661;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27623;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27599;
    wire N__27598;
    wire N__27595;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27565;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27545;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27520;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27505;
    wire N__27500;
    wire N__27497;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27475;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27452;
    wire N__27451;
    wire N__27446;
    wire N__27443;
    wire N__27440;
    wire N__27439;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27394;
    wire N__27391;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27358;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27346;
    wire N__27343;
    wire N__27340;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27321;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27305;
    wire N__27304;
    wire N__27301;
    wire N__27296;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27274;
    wire N__27271;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27244;
    wire N__27239;
    wire N__27238;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27224;
    wire N__27221;
    wire N__27220;
    wire N__27215;
    wire N__27212;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27176;
    wire N__27173;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27121;
    wire N__27120;
    wire N__27117;
    wire N__27116;
    wire N__27115;
    wire N__27114;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27094;
    wire N__27091;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27073;
    wire N__27070;
    wire N__27059;
    wire N__27054;
    wire N__27049;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26947;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26935;
    wire N__26930;
    wire N__26929;
    wire N__26928;
    wire N__26925;
    wire N__26920;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26905;
    wire N__26900;
    wire N__26897;
    wire N__26896;
    wire N__26893;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26842;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26830;
    wire N__26825;
    wire N__26824;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26812;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26794;
    wire N__26789;
    wire N__26786;
    wire N__26785;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26756;
    wire N__26753;
    wire N__26750;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26464;
    wire N__26459;
    wire N__26456;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26444;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26380;
    wire N__26377;
    wire N__26374;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26324;
    wire N__26321;
    wire N__26320;
    wire N__26319;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26303;
    wire N__26300;
    wire N__26299;
    wire N__26298;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26210;
    wire N__26209;
    wire N__26208;
    wire N__26207;
    wire N__26206;
    wire N__26205;
    wire N__26204;
    wire N__26203;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26199;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26195;
    wire N__26194;
    wire N__26193;
    wire N__26192;
    wire N__26189;
    wire N__26182;
    wire N__26181;
    wire N__26180;
    wire N__26179;
    wire N__26178;
    wire N__26177;
    wire N__26176;
    wire N__26175;
    wire N__26174;
    wire N__26173;
    wire N__26172;
    wire N__26171;
    wire N__26170;
    wire N__26169;
    wire N__26162;
    wire N__26153;
    wire N__26144;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26117;
    wire N__26108;
    wire N__26099;
    wire N__26096;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26080;
    wire N__26067;
    wire N__26064;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26041;
    wire N__26040;
    wire N__26037;
    wire N__26032;
    wire N__26027;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25996;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25957;
    wire N__25954;
    wire N__25953;
    wire N__25950;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25928;
    wire N__25925;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25914;
    wire N__25911;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25882;
    wire N__25881;
    wire N__25878;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25708;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25618;
    wire N__25617;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25599;
    wire N__25592;
    wire N__25589;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25567;
    wire N__25564;
    wire N__25563;
    wire N__25560;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25538;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25526;
    wire N__25523;
    wire N__25522;
    wire N__25521;
    wire N__25518;
    wire N__25517;
    wire N__25516;
    wire N__25515;
    wire N__25514;
    wire N__25513;
    wire N__25512;
    wire N__25511;
    wire N__25510;
    wire N__25509;
    wire N__25508;
    wire N__25507;
    wire N__25506;
    wire N__25505;
    wire N__25504;
    wire N__25503;
    wire N__25502;
    wire N__25501;
    wire N__25496;
    wire N__25487;
    wire N__25480;
    wire N__25479;
    wire N__25476;
    wire N__25475;
    wire N__25474;
    wire N__25473;
    wire N__25472;
    wire N__25471;
    wire N__25470;
    wire N__25467;
    wire N__25462;
    wire N__25447;
    wire N__25440;
    wire N__25437;
    wire N__25436;
    wire N__25435;
    wire N__25432;
    wire N__25419;
    wire N__25414;
    wire N__25409;
    wire N__25408;
    wire N__25405;
    wire N__25404;
    wire N__25403;
    wire N__25398;
    wire N__25393;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25358;
    wire N__25355;
    wire N__25354;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25319;
    wire N__25318;
    wire N__25317;
    wire N__25314;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25289;
    wire N__25288;
    wire N__25283;
    wire N__25282;
    wire N__25281;
    wire N__25280;
    wire N__25277;
    wire N__25270;
    wire N__25269;
    wire N__25268;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25243;
    wire N__25242;
    wire N__25241;
    wire N__25240;
    wire N__25237;
    wire N__25236;
    wire N__25235;
    wire N__25228;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25216;
    wire N__25215;
    wire N__25214;
    wire N__25211;
    wire N__25206;
    wire N__25201;
    wire N__25196;
    wire N__25191;
    wire N__25188;
    wire N__25181;
    wire N__25180;
    wire N__25179;
    wire N__25176;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25154;
    wire N__25153;
    wire N__25152;
    wire N__25151;
    wire N__25148;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25140;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25109;
    wire N__25108;
    wire N__25107;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25069;
    wire N__25066;
    wire N__25065;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25038;
    wire N__25031;
    wire N__25030;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25012;
    wire N__25011;
    wire N__25010;
    wire N__25007;
    wire N__25002;
    wire N__24999;
    wire N__24994;
    wire N__24989;
    wire N__24986;
    wire N__24985;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24963;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24943;
    wire N__24938;
    wire N__24937;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24916;
    wire N__24915;
    wire N__24912;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24894;
    wire N__24887;
    wire N__24886;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24865;
    wire N__24864;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24840;
    wire N__24833;
    wire N__24832;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24807;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24795;
    wire N__24788;
    wire N__24787;
    wire N__24784;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24772;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24726;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24695;
    wire N__24694;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24679;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24668;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24641;
    wire N__24640;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24628;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24614;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24593;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24534;
    wire N__24527;
    wire N__24526;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24501;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24470;
    wire N__24469;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24454;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24435;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24419;
    wire N__24418;
    wire N__24415;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24400;
    wire N__24397;
    wire N__24396;
    wire N__24393;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24369;
    wire N__24362;
    wire N__24359;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24337;
    wire N__24334;
    wire N__24333;
    wire N__24330;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24310;
    wire N__24305;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24277;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24256;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24239;
    wire N__24238;
    wire N__24237;
    wire N__24234;
    wire N__24229;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24208;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24158;
    wire N__24157;
    wire N__24156;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24144;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24115;
    wire N__24112;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24081;
    wire N__24078;
    wire N__24071;
    wire N__24070;
    wire N__24067;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24032;
    wire N__24029;
    wire N__24028;
    wire N__24025;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24007;
    wire N__24004;
    wire N__24003;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23974;
    wire N__23973;
    wire N__23970;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23932;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23921;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23903;
    wire N__23902;
    wire N__23901;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23889;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23848;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23838;
    wire N__23835;
    wire N__23834;
    wire N__23829;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23765;
    wire N__23762;
    wire N__23761;
    wire N__23758;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23737;
    wire N__23736;
    wire N__23731;
    wire N__23728;
    wire N__23723;
    wire N__23722;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23678;
    wire N__23675;
    wire N__23674;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23660;
    wire N__23655;
    wire N__23652;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23613;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23476;
    wire N__23475;
    wire N__23474;
    wire N__23473;
    wire N__23472;
    wire N__23471;
    wire N__23470;
    wire N__23469;
    wire N__23468;
    wire N__23467;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23440;
    wire N__23439;
    wire N__23438;
    wire N__23437;
    wire N__23436;
    wire N__23431;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23427;
    wire N__23426;
    wire N__23425;
    wire N__23424;
    wire N__23423;
    wire N__23422;
    wire N__23421;
    wire N__23420;
    wire N__23417;
    wire N__23410;
    wire N__23403;
    wire N__23390;
    wire N__23387;
    wire N__23386;
    wire N__23385;
    wire N__23380;
    wire N__23377;
    wire N__23362;
    wire N__23353;
    wire N__23350;
    wire N__23345;
    wire N__23340;
    wire N__23335;
    wire N__23330;
    wire N__23321;
    wire N__23318;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23284;
    wire N__23283;
    wire N__23282;
    wire N__23281;
    wire N__23280;
    wire N__23279;
    wire N__23278;
    wire N__23277;
    wire N__23276;
    wire N__23275;
    wire N__23274;
    wire N__23273;
    wire N__23272;
    wire N__23271;
    wire N__23270;
    wire N__23269;
    wire N__23268;
    wire N__23265;
    wire N__23264;
    wire N__23263;
    wire N__23262;
    wire N__23259;
    wire N__23258;
    wire N__23245;
    wire N__23240;
    wire N__23233;
    wire N__23226;
    wire N__23225;
    wire N__23224;
    wire N__23223;
    wire N__23222;
    wire N__23221;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23209;
    wire N__23200;
    wire N__23197;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23182;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23150;
    wire N__23145;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23119;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22057;
    wire N__22056;
    wire N__22053;
    wire N__22048;
    wire N__22045;
    wire N__22040;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21837;
    wire N__21834;
    wire N__21829;
    wire N__21826;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21797;
    wire N__21794;
    wire N__21793;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21767;
    wire N__21764;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21745;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21727;
    wire N__21724;
    wire N__21719;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21649;
    wire N__21646;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21592;
    wire N__21591;
    wire N__21590;
    wire N__21589;
    wire N__21588;
    wire N__21587;
    wire N__21586;
    wire N__21585;
    wire N__21584;
    wire N__21573;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21520;
    wire N__21517;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21493;
    wire N__21490;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21475;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21448;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21397;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21358;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21319;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21280;
    wire N__21277;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21238;
    wire N__21235;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21196;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21176;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21164;
    wire N__21161;
    wire N__21160;
    wire N__21159;
    wire N__21156;
    wire N__21151;
    wire N__21146;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21121;
    wire N__21120;
    wire N__21117;
    wire N__21112;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21086;
    wire N__21083;
    wire N__21082;
    wire N__21081;
    wire N__21078;
    wire N__21073;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21055;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21016;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21001;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20977;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20944;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20746;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20713;
    wire N__20710;
    wire N__20709;
    wire N__20708;
    wire N__20707;
    wire N__20704;
    wire N__20703;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20695;
    wire N__20692;
    wire N__20691;
    wire N__20690;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20678;
    wire N__20675;
    wire N__20668;
    wire N__20665;
    wire N__20660;
    wire N__20655;
    wire N__20652;
    wire N__20645;
    wire N__20636;
    wire N__20633;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20564;
    wire N__20563;
    wire N__20562;
    wire N__20561;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20533;
    wire N__20532;
    wire N__20531;
    wire N__20530;
    wire N__20529;
    wire N__20526;
    wire N__20523;
    wire N__20514;
    wire N__20507;
    wire N__20504;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20365;
    wire N__20364;
    wire N__20363;
    wire N__20362;
    wire N__20361;
    wire N__20358;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20346;
    wire N__20345;
    wire N__20344;
    wire N__20343;
    wire N__20340;
    wire N__20339;
    wire N__20338;
    wire N__20337;
    wire N__20336;
    wire N__20335;
    wire N__20334;
    wire N__20333;
    wire N__20332;
    wire N__20331;
    wire N__20330;
    wire N__20329;
    wire N__20328;
    wire N__20327;
    wire N__20326;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20322;
    wire N__20321;
    wire N__20320;
    wire N__20319;
    wire N__20310;
    wire N__20307;
    wire N__20300;
    wire N__20297;
    wire N__20286;
    wire N__20285;
    wire N__20268;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20242;
    wire N__20237;
    wire N__20234;
    wire N__20229;
    wire N__20226;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20207;
    wire N__20198;
    wire N__20195;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20167;
    wire N__20166;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20162;
    wire N__20161;
    wire N__20160;
    wire N__20159;
    wire N__20150;
    wire N__20145;
    wire N__20136;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19809;
    wire N__19808;
    wire N__19807;
    wire N__19802;
    wire N__19801;
    wire N__19798;
    wire N__19797;
    wire N__19794;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19774;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire bfn_1_15_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_1_16_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire bfn_1_17_0_;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire bfn_1_18_0_;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire bfn_1_19_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire bfn_1_20_0_;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire bfn_1_21_0_;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire bfn_1_22_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire bfn_1_23_0_;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire bfn_1_24_0_;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire N_86_i_i;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ;
    wire N_19_1;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_2_21_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_2_22_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire bfn_2_23_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire un7_start_stop;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_3_16_0_;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_3_17_0_;
    wire \pwm_generator_inst.threshold_9 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \pwm_generator_inst.N_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.N_98_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.N_96_cascade_ ;
    wire pwm_duty_input_6;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire pwm_duty_input_3;
    wire pwm_duty_input_5;
    wire pwm_duty_input_7;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire bfn_4_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire bfn_4_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire bfn_4_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire bfn_4_15_0_;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.N_77 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire pwm_duty_input_0;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire pwm_duty_input_1;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire bfn_5_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire bfn_5_15_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.N_46 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire bfn_5_19_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire bfn_5_20_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire bfn_5_21_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire bfn_5_22_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire pwm_duty_input_8;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.N_158 ;
    wire pwm_duty_input_9;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire bfn_7_10_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire bfn_7_11_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_7_12_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_7_13_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.N_160 ;
    wire pwm_duty_input_2;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_8_10_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_8_11_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire bfn_8_12_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8_cascade_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_27 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire elapsed_time_ns_1_RNIT6OBB_0_10_cascade_;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire elapsed_time_ns_1_RNILK91B_0_9_cascade_;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire elapsed_time_ns_1_RNI2COBB_0_15_cascade_;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire elapsed_time_ns_1_RNI5GPBB_0_27_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire s3_phy_c;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_10_9_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_10_10_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire bfn_10_11_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire elapsed_time_ns_1_RNI7IPBB_0_29_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.test_0_sqmuxa ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.N_58 ;
    wire \phase_controller_inst2.N_51_0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_28 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire s4_phy_c;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire elapsed_time_ns_1_RNI4EOBB_0_17_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.N_49_0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire bfn_11_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_11_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_11_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_11_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire start_stop_c;
    wire il_max_comp2_c;
    wire phase_controller_inst1_N_54_cascade_;
    wire \phase_controller_inst2.N_54 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.N_166_i ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_11_19_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire bfn_11_20_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire bfn_11_21_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire bfn_11_22_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_27 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_28 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_30 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_31 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire test22_c;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire bfn_12_10_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_12_11_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_12_12_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_12_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \phase_controller_inst1.N_52 ;
    wire phase_controller_inst1_N_54;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.N_1271_i ;
    wire \current_shift_inst.control_input_1 ;
    wire bfn_12_17_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_12_18_0_;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.control_input_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire \current_shift_inst.control_input_cry_14 ;
    wire \current_shift_inst.control_input_cry_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire bfn_12_19_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.control_input_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.control_input_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.control_input_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.control_input_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.control_input_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.control_input_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.control_input_cry_22 ;
    wire \current_shift_inst.control_input_cry_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire bfn_12_20_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.control_input_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ;
    wire \current_shift_inst.control_input_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ;
    wire \current_shift_inst.control_input_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ;
    wire \current_shift_inst.control_input_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ;
    wire \current_shift_inst.control_input_cry_28 ;
    wire \current_shift_inst.control_input_cry_29 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ;
    wire \pll_inst.red_c_i ;
    wire il_min_comp1_c;
    wire \phase_controller_inst1.N_56 ;
    wire phase_controller_inst1_state_4;
    wire elapsed_time_ns_1_RNIH33T9_0_5_cascade_;
    wire elapsed_time_ns_1_RNIU0DN9_0_20_cascade_;
    wire \phase_controller_inst1.test_0_sqmuxa ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire bfn_13_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire bfn_13_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire bfn_13_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_13_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_165_i ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire il_max_comp1_c;
    wire test_c;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.control_input_axb_16 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.control_input_axb_18 ;
    wire \current_shift_inst.control_input_axb_17 ;
    wire \current_shift_inst.control_input_axb_20 ;
    wire \current_shift_inst.control_input_axb_21 ;
    wire \current_shift_inst.control_input_axb_22 ;
    wire \current_shift_inst.control_input_axb_27 ;
    wire \current_shift_inst.control_input_axb_26 ;
    wire \current_shift_inst.control_input_axb_25 ;
    wire \current_shift_inst.control_input_axb_29 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire s1_phy_c;
    wire state_3;
    wire \current_shift_inst.timer_s1.N_161_i ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire delay_hc_input_c_g;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_14_4_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_14_5_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire bfn_14_6_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire bfn_14_10_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_14_11_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_14_12_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_14_13_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ;
    wire \current_shift_inst.un38_control_input_0_s0_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.control_input_axb_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_15_5_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_15_6_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_15_7_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_15_8_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_15_10_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_15_11_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire bfn_15_12_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire bfn_15_13_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ;
    wire \current_shift_inst.un38_control_input_0_s1_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire bfn_15_14_0_;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_15_15_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_15_16_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.control_input_axb_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire \current_shift_inst.control_input_axb_13 ;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.control_input_axb_14 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.control_input_axb_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.control_input_axb_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire bfn_16_17_0_;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_16_18_0_;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_16_19_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_16_20_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire elapsed_time_ns_1_RNI46CN9_0_17_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire elapsed_time_ns_1_RNITUBN9_0_10_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire elapsed_time_ns_1_RNI02CN9_0_13_cascade_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_17_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_17_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.N_164_i ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire bfn_17_15_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_17_16_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_17_17_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire bfn_18_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_18_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire bfn_18_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_18_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.N_163_i ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_18_19_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_18_20_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_18_21_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire bfn_18_22_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_161_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_18_23_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_18_24_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_18_25_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_18_26_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_162_i ;
    wire GB_BUFFER_clock_output_0_THRU_CO;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire _gnd_net_;
    wire clock_output_0;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__27917),
            .RESETB(N__33224),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clock_output_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__44835),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__44832),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__30764,N__30791,N__30821,N__30848,N__30881,N__30911,N__30941,N__30971,N__30512,N__30542,N__30569,N__30599,N__30632,N__30662,N__30698,N__30728}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__44834,dangling_wire_45,N__44833}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__44965),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__44891),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__20333,N__20326,N__20331,N__20325,N__20332,N__20324,N__20334,N__20321,N__20327,N__20320,N__20328,N__20322,N__20329,N__20323,N__20330}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__44964,N__44894,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__44892,N__44963,N__44893,N__44962}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__44715),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__44708),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__20343,N__20362,N__20344,N__20363,N__20345,N__25107,N__25319,N__22061,N__21845,N__21718,N__21792,N__21746,N__26026,N__22559,N__22589}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__44714,N__44711,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__44709,N__44713,N__44710,N__44712}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__44816),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__44813),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__30242,N__30275,N__30299,N__30329,N__30359,N__30389,N__30422,N__30448,N__30488,N__30071,N__30107,N__30137,N__30170,N__30206,N__29636}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__44815,dangling_wire_215,N__44814}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__51009),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__51011),
            .DIN(N__51010),
            .DOUT(N__51009),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__51011),
            .PADOUT(N__51010),
            .PADIN(N__51009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clock_output_obuf_iopad (
            .OE(N__51000),
            .DIN(N__50999),
            .DOUT(N__50998),
            .PACKAGEPIN(clock_output));
    defparam clock_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam clock_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO clock_output_obuf_preio (
            .PADOEN(N__51000),
            .PADOUT(N__50999),
            .PADIN(N__50998),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__50597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test_obuf_iopad (
            .OE(N__50991),
            .DIN(N__50990),
            .DOUT(N__50989),
            .PACKAGEPIN(test));
    defparam test_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test_obuf_preio (
            .PADOEN(N__50991),
            .PADOUT(N__50990),
            .PADIN(N__50989),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35621),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__50982),
            .DIN(N__50981),
            .DOUT(N__50980),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__50982),
            .PADOUT(N__50981),
            .PADIN(N__50980),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__50973),
            .DIN(N__50972),
            .DOUT(N__50971),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__50973),
            .PADOUT(N__50972),
            .PADIN(N__50971),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__50964),
            .DIN(N__50963),
            .DOUT(N__50962),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__50964),
            .PADOUT(N__50963),
            .PADIN(N__50962),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21620),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__50955),
            .DIN(N__50954),
            .DOUT(N__50953),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__50955),
            .PADOUT(N__50954),
            .PADIN(N__50953),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__50946),
            .DIN(N__50945),
            .DOUT(N__50944),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__50946),
            .PADOUT(N__50945),
            .PADIN(N__50944),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35774),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test22_obuf_iopad (
            .OE(N__50937),
            .DIN(N__50936),
            .DOUT(N__50935),
            .PACKAGEPIN(test22));
    defparam test22_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test22_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test22_obuf_preio (
            .PADOEN(N__50937),
            .PADOUT(N__50936),
            .PADIN(N__50935),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31007),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__50928),
            .DIN(N__50927),
            .DOUT(N__50926),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__50928),
            .PADOUT(N__50927),
            .PADIN(N__50926),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__50919),
            .DIN(N__50918),
            .DOUT(N__50917),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__50919),
            .PADOUT(N__50918),
            .PADIN(N__50917),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35924),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__50910),
            .DIN(N__50909),
            .DOUT(N__50908),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__50910),
            .PADOUT(N__50909),
            .PADIN(N__50908),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28994),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__50901),
            .DIN(N__50900),
            .DOUT(N__50899),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__50901),
            .PADOUT(N__50900),
            .PADIN(N__50899),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__50892),
            .DIN(N__50891),
            .DOUT(N__50890),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__50892),
            .PADOUT(N__50891),
            .PADIN(N__50890),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27938),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__50883),
            .DIN(N__50882),
            .DOUT(N__50881),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__50883),
            .PADOUT(N__50882),
            .PADIN(N__50881),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__50874),
            .DIN(N__50873),
            .DOUT(N__50872),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__50874),
            .PADOUT(N__50873),
            .PADIN(N__50872),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__12164 (
            .O(N__50855),
            .I(N__50852));
    InMux I__12163 (
            .O(N__50852),
            .I(N__50847));
    InMux I__12162 (
            .O(N__50851),
            .I(N__50844));
    InMux I__12161 (
            .O(N__50850),
            .I(N__50841));
    LocalMux I__12160 (
            .O(N__50847),
            .I(N__50836));
    LocalMux I__12159 (
            .O(N__50844),
            .I(N__50836));
    LocalMux I__12158 (
            .O(N__50841),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv12 I__12157 (
            .O(N__50836),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__12156 (
            .O(N__50831),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__12155 (
            .O(N__50828),
            .I(N__50824));
    CascadeMux I__12154 (
            .O(N__50827),
            .I(N__50821));
    InMux I__12153 (
            .O(N__50824),
            .I(N__50815));
    InMux I__12152 (
            .O(N__50821),
            .I(N__50815));
    InMux I__12151 (
            .O(N__50820),
            .I(N__50812));
    LocalMux I__12150 (
            .O(N__50815),
            .I(N__50809));
    LocalMux I__12149 (
            .O(N__50812),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv12 I__12148 (
            .O(N__50809),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__12147 (
            .O(N__50804),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__12146 (
            .O(N__50801),
            .I(N__50797));
    InMux I__12145 (
            .O(N__50800),
            .I(N__50794));
    LocalMux I__12144 (
            .O(N__50797),
            .I(N__50791));
    LocalMux I__12143 (
            .O(N__50794),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv12 I__12142 (
            .O(N__50791),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__12141 (
            .O(N__50786),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__12140 (
            .O(N__50783),
            .I(N__50745));
    InMux I__12139 (
            .O(N__50782),
            .I(N__50745));
    InMux I__12138 (
            .O(N__50781),
            .I(N__50745));
    InMux I__12137 (
            .O(N__50780),
            .I(N__50745));
    InMux I__12136 (
            .O(N__50779),
            .I(N__50736));
    InMux I__12135 (
            .O(N__50778),
            .I(N__50736));
    InMux I__12134 (
            .O(N__50777),
            .I(N__50736));
    InMux I__12133 (
            .O(N__50776),
            .I(N__50736));
    InMux I__12132 (
            .O(N__50775),
            .I(N__50731));
    InMux I__12131 (
            .O(N__50774),
            .I(N__50731));
    InMux I__12130 (
            .O(N__50773),
            .I(N__50722));
    InMux I__12129 (
            .O(N__50772),
            .I(N__50722));
    InMux I__12128 (
            .O(N__50771),
            .I(N__50722));
    InMux I__12127 (
            .O(N__50770),
            .I(N__50722));
    InMux I__12126 (
            .O(N__50769),
            .I(N__50713));
    InMux I__12125 (
            .O(N__50768),
            .I(N__50713));
    InMux I__12124 (
            .O(N__50767),
            .I(N__50713));
    InMux I__12123 (
            .O(N__50766),
            .I(N__50713));
    InMux I__12122 (
            .O(N__50765),
            .I(N__50704));
    InMux I__12121 (
            .O(N__50764),
            .I(N__50704));
    InMux I__12120 (
            .O(N__50763),
            .I(N__50704));
    InMux I__12119 (
            .O(N__50762),
            .I(N__50704));
    InMux I__12118 (
            .O(N__50761),
            .I(N__50695));
    InMux I__12117 (
            .O(N__50760),
            .I(N__50695));
    InMux I__12116 (
            .O(N__50759),
            .I(N__50695));
    InMux I__12115 (
            .O(N__50758),
            .I(N__50695));
    InMux I__12114 (
            .O(N__50757),
            .I(N__50686));
    InMux I__12113 (
            .O(N__50756),
            .I(N__50686));
    InMux I__12112 (
            .O(N__50755),
            .I(N__50686));
    InMux I__12111 (
            .O(N__50754),
            .I(N__50686));
    LocalMux I__12110 (
            .O(N__50745),
            .I(N__50673));
    LocalMux I__12109 (
            .O(N__50736),
            .I(N__50673));
    LocalMux I__12108 (
            .O(N__50731),
            .I(N__50673));
    LocalMux I__12107 (
            .O(N__50722),
            .I(N__50673));
    LocalMux I__12106 (
            .O(N__50713),
            .I(N__50673));
    LocalMux I__12105 (
            .O(N__50704),
            .I(N__50673));
    LocalMux I__12104 (
            .O(N__50695),
            .I(N__50668));
    LocalMux I__12103 (
            .O(N__50686),
            .I(N__50668));
    Span4Mux_v I__12102 (
            .O(N__50673),
            .I(N__50665));
    Odrv12 I__12101 (
            .O(N__50668),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__12100 (
            .O(N__50665),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__12099 (
            .O(N__50660),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__12098 (
            .O(N__50657),
            .I(N__50653));
    InMux I__12097 (
            .O(N__50656),
            .I(N__50650));
    LocalMux I__12096 (
            .O(N__50653),
            .I(N__50647));
    LocalMux I__12095 (
            .O(N__50650),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv12 I__12094 (
            .O(N__50647),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__12093 (
            .O(N__50642),
            .I(N__50637));
    CEMux I__12092 (
            .O(N__50641),
            .I(N__50634));
    CEMux I__12091 (
            .O(N__50640),
            .I(N__50630));
    LocalMux I__12090 (
            .O(N__50637),
            .I(N__50625));
    LocalMux I__12089 (
            .O(N__50634),
            .I(N__50625));
    CEMux I__12088 (
            .O(N__50633),
            .I(N__50622));
    LocalMux I__12087 (
            .O(N__50630),
            .I(N__50619));
    Span4Mux_v I__12086 (
            .O(N__50625),
            .I(N__50616));
    LocalMux I__12085 (
            .O(N__50622),
            .I(N__50613));
    Span4Mux_h I__12084 (
            .O(N__50619),
            .I(N__50610));
    Span4Mux_h I__12083 (
            .O(N__50616),
            .I(N__50607));
    Span4Mux_h I__12082 (
            .O(N__50613),
            .I(N__50604));
    Odrv4 I__12081 (
            .O(N__50610),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    Odrv4 I__12080 (
            .O(N__50607),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    Odrv4 I__12079 (
            .O(N__50604),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    IoInMux I__12078 (
            .O(N__50597),
            .I(N__50594));
    LocalMux I__12077 (
            .O(N__50594),
            .I(GB_BUFFER_clock_output_0_THRU_CO));
    InMux I__12076 (
            .O(N__50591),
            .I(N__50585));
    InMux I__12075 (
            .O(N__50590),
            .I(N__50580));
    InMux I__12074 (
            .O(N__50589),
            .I(N__50580));
    InMux I__12073 (
            .O(N__50588),
            .I(N__50577));
    LocalMux I__12072 (
            .O(N__50585),
            .I(N__50574));
    LocalMux I__12071 (
            .O(N__50580),
            .I(N__50571));
    LocalMux I__12070 (
            .O(N__50577),
            .I(N__50568));
    Span4Mux_v I__12069 (
            .O(N__50574),
            .I(N__50563));
    Span4Mux_v I__12068 (
            .O(N__50571),
            .I(N__50563));
    Odrv4 I__12067 (
            .O(N__50568),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__12066 (
            .O(N__50563),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__12065 (
            .O(N__50558),
            .I(N__50553));
    InMux I__12064 (
            .O(N__50557),
            .I(N__50550));
    InMux I__12063 (
            .O(N__50556),
            .I(N__50547));
    LocalMux I__12062 (
            .O(N__50553),
            .I(N__50544));
    LocalMux I__12061 (
            .O(N__50550),
            .I(N__50541));
    LocalMux I__12060 (
            .O(N__50547),
            .I(N__50536));
    Span4Mux_v I__12059 (
            .O(N__50544),
            .I(N__50536));
    Span12Mux_s9_h I__12058 (
            .O(N__50541),
            .I(N__50533));
    Odrv4 I__12057 (
            .O(N__50536),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv12 I__12056 (
            .O(N__50533),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__12055 (
            .O(N__50528),
            .I(N__50502));
    InMux I__12054 (
            .O(N__50527),
            .I(N__50490));
    InMux I__12053 (
            .O(N__50526),
            .I(N__50487));
    CascadeMux I__12052 (
            .O(N__50525),
            .I(N__50474));
    InMux I__12051 (
            .O(N__50524),
            .I(N__50470));
    InMux I__12050 (
            .O(N__50523),
            .I(N__50464));
    InMux I__12049 (
            .O(N__50522),
            .I(N__50464));
    InMux I__12048 (
            .O(N__50521),
            .I(N__50461));
    InMux I__12047 (
            .O(N__50520),
            .I(N__50458));
    InMux I__12046 (
            .O(N__50519),
            .I(N__50449));
    InMux I__12045 (
            .O(N__50518),
            .I(N__50449));
    InMux I__12044 (
            .O(N__50517),
            .I(N__50449));
    InMux I__12043 (
            .O(N__50516),
            .I(N__50449));
    InMux I__12042 (
            .O(N__50515),
            .I(N__50442));
    InMux I__12041 (
            .O(N__50514),
            .I(N__50442));
    InMux I__12040 (
            .O(N__50513),
            .I(N__50442));
    InMux I__12039 (
            .O(N__50512),
            .I(N__50435));
    InMux I__12038 (
            .O(N__50511),
            .I(N__50435));
    InMux I__12037 (
            .O(N__50510),
            .I(N__50435));
    InMux I__12036 (
            .O(N__50509),
            .I(N__50424));
    InMux I__12035 (
            .O(N__50508),
            .I(N__50424));
    InMux I__12034 (
            .O(N__50507),
            .I(N__50424));
    InMux I__12033 (
            .O(N__50506),
            .I(N__50424));
    InMux I__12032 (
            .O(N__50505),
            .I(N__50424));
    LocalMux I__12031 (
            .O(N__50502),
            .I(N__50421));
    InMux I__12030 (
            .O(N__50501),
            .I(N__50417));
    InMux I__12029 (
            .O(N__50500),
            .I(N__50412));
    InMux I__12028 (
            .O(N__50499),
            .I(N__50412));
    CascadeMux I__12027 (
            .O(N__50498),
            .I(N__50391));
    InMux I__12026 (
            .O(N__50497),
            .I(N__50381));
    InMux I__12025 (
            .O(N__50496),
            .I(N__50381));
    InMux I__12024 (
            .O(N__50495),
            .I(N__50381));
    InMux I__12023 (
            .O(N__50494),
            .I(N__50381));
    InMux I__12022 (
            .O(N__50493),
            .I(N__50378));
    LocalMux I__12021 (
            .O(N__50490),
            .I(N__50375));
    LocalMux I__12020 (
            .O(N__50487),
            .I(N__50372));
    InMux I__12019 (
            .O(N__50486),
            .I(N__50367));
    InMux I__12018 (
            .O(N__50485),
            .I(N__50367));
    InMux I__12017 (
            .O(N__50484),
            .I(N__50364));
    InMux I__12016 (
            .O(N__50483),
            .I(N__50355));
    InMux I__12015 (
            .O(N__50482),
            .I(N__50355));
    InMux I__12014 (
            .O(N__50481),
            .I(N__50355));
    InMux I__12013 (
            .O(N__50480),
            .I(N__50355));
    InMux I__12012 (
            .O(N__50479),
            .I(N__50340));
    InMux I__12011 (
            .O(N__50478),
            .I(N__50340));
    InMux I__12010 (
            .O(N__50477),
            .I(N__50340));
    InMux I__12009 (
            .O(N__50474),
            .I(N__50340));
    InMux I__12008 (
            .O(N__50473),
            .I(N__50340));
    LocalMux I__12007 (
            .O(N__50470),
            .I(N__50337));
    InMux I__12006 (
            .O(N__50469),
            .I(N__50334));
    LocalMux I__12005 (
            .O(N__50464),
            .I(N__50322));
    LocalMux I__12004 (
            .O(N__50461),
            .I(N__50319));
    LocalMux I__12003 (
            .O(N__50458),
            .I(N__50314));
    LocalMux I__12002 (
            .O(N__50449),
            .I(N__50314));
    LocalMux I__12001 (
            .O(N__50442),
            .I(N__50311));
    LocalMux I__12000 (
            .O(N__50435),
            .I(N__50304));
    LocalMux I__11999 (
            .O(N__50424),
            .I(N__50304));
    Span4Mux_h I__11998 (
            .O(N__50421),
            .I(N__50304));
    CascadeMux I__11997 (
            .O(N__50420),
            .I(N__50299));
    LocalMux I__11996 (
            .O(N__50417),
            .I(N__50287));
    LocalMux I__11995 (
            .O(N__50412),
            .I(N__50284));
    InMux I__11994 (
            .O(N__50411),
            .I(N__50276));
    InMux I__11993 (
            .O(N__50410),
            .I(N__50276));
    InMux I__11992 (
            .O(N__50409),
            .I(N__50265));
    InMux I__11991 (
            .O(N__50408),
            .I(N__50265));
    InMux I__11990 (
            .O(N__50407),
            .I(N__50265));
    InMux I__11989 (
            .O(N__50406),
            .I(N__50265));
    InMux I__11988 (
            .O(N__50405),
            .I(N__50265));
    InMux I__11987 (
            .O(N__50404),
            .I(N__50256));
    InMux I__11986 (
            .O(N__50403),
            .I(N__50256));
    InMux I__11985 (
            .O(N__50402),
            .I(N__50256));
    InMux I__11984 (
            .O(N__50401),
            .I(N__50256));
    InMux I__11983 (
            .O(N__50400),
            .I(N__50251));
    InMux I__11982 (
            .O(N__50399),
            .I(N__50251));
    InMux I__11981 (
            .O(N__50398),
            .I(N__50248));
    InMux I__11980 (
            .O(N__50397),
            .I(N__50245));
    InMux I__11979 (
            .O(N__50396),
            .I(N__50234));
    InMux I__11978 (
            .O(N__50395),
            .I(N__50234));
    InMux I__11977 (
            .O(N__50394),
            .I(N__50234));
    InMux I__11976 (
            .O(N__50391),
            .I(N__50234));
    InMux I__11975 (
            .O(N__50390),
            .I(N__50234));
    LocalMux I__11974 (
            .O(N__50381),
            .I(N__50219));
    LocalMux I__11973 (
            .O(N__50378),
            .I(N__50219));
    Span4Mux_s3_v I__11972 (
            .O(N__50375),
            .I(N__50219));
    Span4Mux_v I__11971 (
            .O(N__50372),
            .I(N__50219));
    LocalMux I__11970 (
            .O(N__50367),
            .I(N__50219));
    LocalMux I__11969 (
            .O(N__50364),
            .I(N__50219));
    LocalMux I__11968 (
            .O(N__50355),
            .I(N__50219));
    InMux I__11967 (
            .O(N__50354),
            .I(N__50210));
    InMux I__11966 (
            .O(N__50353),
            .I(N__50210));
    InMux I__11965 (
            .O(N__50352),
            .I(N__50210));
    InMux I__11964 (
            .O(N__50351),
            .I(N__50210));
    LocalMux I__11963 (
            .O(N__50340),
            .I(N__50207));
    Span4Mux_v I__11962 (
            .O(N__50337),
            .I(N__50202));
    LocalMux I__11961 (
            .O(N__50334),
            .I(N__50202));
    InMux I__11960 (
            .O(N__50333),
            .I(N__50189));
    InMux I__11959 (
            .O(N__50332),
            .I(N__50189));
    InMux I__11958 (
            .O(N__50331),
            .I(N__50189));
    InMux I__11957 (
            .O(N__50330),
            .I(N__50189));
    InMux I__11956 (
            .O(N__50329),
            .I(N__50189));
    InMux I__11955 (
            .O(N__50328),
            .I(N__50189));
    InMux I__11954 (
            .O(N__50327),
            .I(N__50182));
    InMux I__11953 (
            .O(N__50326),
            .I(N__50182));
    InMux I__11952 (
            .O(N__50325),
            .I(N__50182));
    Span4Mux_h I__11951 (
            .O(N__50322),
            .I(N__50173));
    Span4Mux_v I__11950 (
            .O(N__50319),
            .I(N__50173));
    Span4Mux_v I__11949 (
            .O(N__50314),
            .I(N__50173));
    Span4Mux_v I__11948 (
            .O(N__50311),
            .I(N__50173));
    Span4Mux_v I__11947 (
            .O(N__50304),
            .I(N__50170));
    InMux I__11946 (
            .O(N__50303),
            .I(N__50165));
    InMux I__11945 (
            .O(N__50302),
            .I(N__50165));
    InMux I__11944 (
            .O(N__50299),
            .I(N__50160));
    InMux I__11943 (
            .O(N__50298),
            .I(N__50160));
    InMux I__11942 (
            .O(N__50297),
            .I(N__50151));
    InMux I__11941 (
            .O(N__50296),
            .I(N__50151));
    InMux I__11940 (
            .O(N__50295),
            .I(N__50151));
    InMux I__11939 (
            .O(N__50294),
            .I(N__50151));
    InMux I__11938 (
            .O(N__50293),
            .I(N__50142));
    InMux I__11937 (
            .O(N__50292),
            .I(N__50142));
    InMux I__11936 (
            .O(N__50291),
            .I(N__50142));
    InMux I__11935 (
            .O(N__50290),
            .I(N__50142));
    Span4Mux_v I__11934 (
            .O(N__50287),
            .I(N__50137));
    Span4Mux_h I__11933 (
            .O(N__50284),
            .I(N__50137));
    InMux I__11932 (
            .O(N__50283),
            .I(N__50130));
    InMux I__11931 (
            .O(N__50282),
            .I(N__50130));
    InMux I__11930 (
            .O(N__50281),
            .I(N__50130));
    LocalMux I__11929 (
            .O(N__50276),
            .I(N__50123));
    LocalMux I__11928 (
            .O(N__50265),
            .I(N__50123));
    LocalMux I__11927 (
            .O(N__50256),
            .I(N__50123));
    LocalMux I__11926 (
            .O(N__50251),
            .I(N__50116));
    LocalMux I__11925 (
            .O(N__50248),
            .I(N__50116));
    LocalMux I__11924 (
            .O(N__50245),
            .I(N__50116));
    LocalMux I__11923 (
            .O(N__50234),
            .I(N__50111));
    Span4Mux_v I__11922 (
            .O(N__50219),
            .I(N__50111));
    LocalMux I__11921 (
            .O(N__50210),
            .I(N__50104));
    Span4Mux_v I__11920 (
            .O(N__50207),
            .I(N__50104));
    Span4Mux_h I__11919 (
            .O(N__50202),
            .I(N__50104));
    LocalMux I__11918 (
            .O(N__50189),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11917 (
            .O(N__50182),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11916 (
            .O(N__50173),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11915 (
            .O(N__50170),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11914 (
            .O(N__50165),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11913 (
            .O(N__50160),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11912 (
            .O(N__50151),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11911 (
            .O(N__50142),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11910 (
            .O(N__50137),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__11909 (
            .O(N__50130),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11908 (
            .O(N__50123),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__11907 (
            .O(N__50116),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11906 (
            .O(N__50111),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11905 (
            .O(N__50104),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    CascadeMux I__11904 (
            .O(N__50075),
            .I(N__50071));
    CascadeMux I__11903 (
            .O(N__50074),
            .I(N__50068));
    InMux I__11902 (
            .O(N__50071),
            .I(N__50063));
    InMux I__11901 (
            .O(N__50068),
            .I(N__50063));
    LocalMux I__11900 (
            .O(N__50063),
            .I(N__50060));
    Span4Mux_h I__11899 (
            .O(N__50060),
            .I(N__50057));
    Odrv4 I__11898 (
            .O(N__50057),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    InMux I__11897 (
            .O(N__50054),
            .I(N__50051));
    LocalMux I__11896 (
            .O(N__50051),
            .I(N__49896));
    ClkMux I__11895 (
            .O(N__50050),
            .I(N__49583));
    ClkMux I__11894 (
            .O(N__50049),
            .I(N__49583));
    ClkMux I__11893 (
            .O(N__50048),
            .I(N__49583));
    ClkMux I__11892 (
            .O(N__50047),
            .I(N__49583));
    ClkMux I__11891 (
            .O(N__50046),
            .I(N__49583));
    ClkMux I__11890 (
            .O(N__50045),
            .I(N__49583));
    ClkMux I__11889 (
            .O(N__50044),
            .I(N__49583));
    ClkMux I__11888 (
            .O(N__50043),
            .I(N__49583));
    ClkMux I__11887 (
            .O(N__50042),
            .I(N__49583));
    ClkMux I__11886 (
            .O(N__50041),
            .I(N__49583));
    ClkMux I__11885 (
            .O(N__50040),
            .I(N__49583));
    ClkMux I__11884 (
            .O(N__50039),
            .I(N__49583));
    ClkMux I__11883 (
            .O(N__50038),
            .I(N__49583));
    ClkMux I__11882 (
            .O(N__50037),
            .I(N__49583));
    ClkMux I__11881 (
            .O(N__50036),
            .I(N__49583));
    ClkMux I__11880 (
            .O(N__50035),
            .I(N__49583));
    ClkMux I__11879 (
            .O(N__50034),
            .I(N__49583));
    ClkMux I__11878 (
            .O(N__50033),
            .I(N__49583));
    ClkMux I__11877 (
            .O(N__50032),
            .I(N__49583));
    ClkMux I__11876 (
            .O(N__50031),
            .I(N__49583));
    ClkMux I__11875 (
            .O(N__50030),
            .I(N__49583));
    ClkMux I__11874 (
            .O(N__50029),
            .I(N__49583));
    ClkMux I__11873 (
            .O(N__50028),
            .I(N__49583));
    ClkMux I__11872 (
            .O(N__50027),
            .I(N__49583));
    ClkMux I__11871 (
            .O(N__50026),
            .I(N__49583));
    ClkMux I__11870 (
            .O(N__50025),
            .I(N__49583));
    ClkMux I__11869 (
            .O(N__50024),
            .I(N__49583));
    ClkMux I__11868 (
            .O(N__50023),
            .I(N__49583));
    ClkMux I__11867 (
            .O(N__50022),
            .I(N__49583));
    ClkMux I__11866 (
            .O(N__50021),
            .I(N__49583));
    ClkMux I__11865 (
            .O(N__50020),
            .I(N__49583));
    ClkMux I__11864 (
            .O(N__50019),
            .I(N__49583));
    ClkMux I__11863 (
            .O(N__50018),
            .I(N__49583));
    ClkMux I__11862 (
            .O(N__50017),
            .I(N__49583));
    ClkMux I__11861 (
            .O(N__50016),
            .I(N__49583));
    ClkMux I__11860 (
            .O(N__50015),
            .I(N__49583));
    ClkMux I__11859 (
            .O(N__50014),
            .I(N__49583));
    ClkMux I__11858 (
            .O(N__50013),
            .I(N__49583));
    ClkMux I__11857 (
            .O(N__50012),
            .I(N__49583));
    ClkMux I__11856 (
            .O(N__50011),
            .I(N__49583));
    ClkMux I__11855 (
            .O(N__50010),
            .I(N__49583));
    ClkMux I__11854 (
            .O(N__50009),
            .I(N__49583));
    ClkMux I__11853 (
            .O(N__50008),
            .I(N__49583));
    ClkMux I__11852 (
            .O(N__50007),
            .I(N__49583));
    ClkMux I__11851 (
            .O(N__50006),
            .I(N__49583));
    ClkMux I__11850 (
            .O(N__50005),
            .I(N__49583));
    ClkMux I__11849 (
            .O(N__50004),
            .I(N__49583));
    ClkMux I__11848 (
            .O(N__50003),
            .I(N__49583));
    ClkMux I__11847 (
            .O(N__50002),
            .I(N__49583));
    ClkMux I__11846 (
            .O(N__50001),
            .I(N__49583));
    ClkMux I__11845 (
            .O(N__50000),
            .I(N__49583));
    ClkMux I__11844 (
            .O(N__49999),
            .I(N__49583));
    ClkMux I__11843 (
            .O(N__49998),
            .I(N__49583));
    ClkMux I__11842 (
            .O(N__49997),
            .I(N__49583));
    ClkMux I__11841 (
            .O(N__49996),
            .I(N__49583));
    ClkMux I__11840 (
            .O(N__49995),
            .I(N__49583));
    ClkMux I__11839 (
            .O(N__49994),
            .I(N__49583));
    ClkMux I__11838 (
            .O(N__49993),
            .I(N__49583));
    ClkMux I__11837 (
            .O(N__49992),
            .I(N__49583));
    ClkMux I__11836 (
            .O(N__49991),
            .I(N__49583));
    ClkMux I__11835 (
            .O(N__49990),
            .I(N__49583));
    ClkMux I__11834 (
            .O(N__49989),
            .I(N__49583));
    ClkMux I__11833 (
            .O(N__49988),
            .I(N__49583));
    ClkMux I__11832 (
            .O(N__49987),
            .I(N__49583));
    ClkMux I__11831 (
            .O(N__49986),
            .I(N__49583));
    ClkMux I__11830 (
            .O(N__49985),
            .I(N__49583));
    ClkMux I__11829 (
            .O(N__49984),
            .I(N__49583));
    ClkMux I__11828 (
            .O(N__49983),
            .I(N__49583));
    ClkMux I__11827 (
            .O(N__49982),
            .I(N__49583));
    ClkMux I__11826 (
            .O(N__49981),
            .I(N__49583));
    ClkMux I__11825 (
            .O(N__49980),
            .I(N__49583));
    ClkMux I__11824 (
            .O(N__49979),
            .I(N__49583));
    ClkMux I__11823 (
            .O(N__49978),
            .I(N__49583));
    ClkMux I__11822 (
            .O(N__49977),
            .I(N__49583));
    ClkMux I__11821 (
            .O(N__49976),
            .I(N__49583));
    ClkMux I__11820 (
            .O(N__49975),
            .I(N__49583));
    ClkMux I__11819 (
            .O(N__49974),
            .I(N__49583));
    ClkMux I__11818 (
            .O(N__49973),
            .I(N__49583));
    ClkMux I__11817 (
            .O(N__49972),
            .I(N__49583));
    ClkMux I__11816 (
            .O(N__49971),
            .I(N__49583));
    ClkMux I__11815 (
            .O(N__49970),
            .I(N__49583));
    ClkMux I__11814 (
            .O(N__49969),
            .I(N__49583));
    ClkMux I__11813 (
            .O(N__49968),
            .I(N__49583));
    ClkMux I__11812 (
            .O(N__49967),
            .I(N__49583));
    ClkMux I__11811 (
            .O(N__49966),
            .I(N__49583));
    ClkMux I__11810 (
            .O(N__49965),
            .I(N__49583));
    ClkMux I__11809 (
            .O(N__49964),
            .I(N__49583));
    ClkMux I__11808 (
            .O(N__49963),
            .I(N__49583));
    ClkMux I__11807 (
            .O(N__49962),
            .I(N__49583));
    ClkMux I__11806 (
            .O(N__49961),
            .I(N__49583));
    ClkMux I__11805 (
            .O(N__49960),
            .I(N__49583));
    ClkMux I__11804 (
            .O(N__49959),
            .I(N__49583));
    ClkMux I__11803 (
            .O(N__49958),
            .I(N__49583));
    ClkMux I__11802 (
            .O(N__49957),
            .I(N__49583));
    ClkMux I__11801 (
            .O(N__49956),
            .I(N__49583));
    ClkMux I__11800 (
            .O(N__49955),
            .I(N__49583));
    ClkMux I__11799 (
            .O(N__49954),
            .I(N__49583));
    ClkMux I__11798 (
            .O(N__49953),
            .I(N__49583));
    ClkMux I__11797 (
            .O(N__49952),
            .I(N__49583));
    ClkMux I__11796 (
            .O(N__49951),
            .I(N__49583));
    ClkMux I__11795 (
            .O(N__49950),
            .I(N__49583));
    ClkMux I__11794 (
            .O(N__49949),
            .I(N__49583));
    ClkMux I__11793 (
            .O(N__49948),
            .I(N__49583));
    ClkMux I__11792 (
            .O(N__49947),
            .I(N__49583));
    ClkMux I__11791 (
            .O(N__49946),
            .I(N__49583));
    ClkMux I__11790 (
            .O(N__49945),
            .I(N__49583));
    ClkMux I__11789 (
            .O(N__49944),
            .I(N__49583));
    ClkMux I__11788 (
            .O(N__49943),
            .I(N__49583));
    ClkMux I__11787 (
            .O(N__49942),
            .I(N__49583));
    ClkMux I__11786 (
            .O(N__49941),
            .I(N__49583));
    ClkMux I__11785 (
            .O(N__49940),
            .I(N__49583));
    ClkMux I__11784 (
            .O(N__49939),
            .I(N__49583));
    ClkMux I__11783 (
            .O(N__49938),
            .I(N__49583));
    ClkMux I__11782 (
            .O(N__49937),
            .I(N__49583));
    ClkMux I__11781 (
            .O(N__49936),
            .I(N__49583));
    ClkMux I__11780 (
            .O(N__49935),
            .I(N__49583));
    ClkMux I__11779 (
            .O(N__49934),
            .I(N__49583));
    ClkMux I__11778 (
            .O(N__49933),
            .I(N__49583));
    ClkMux I__11777 (
            .O(N__49932),
            .I(N__49583));
    ClkMux I__11776 (
            .O(N__49931),
            .I(N__49583));
    ClkMux I__11775 (
            .O(N__49930),
            .I(N__49583));
    ClkMux I__11774 (
            .O(N__49929),
            .I(N__49583));
    ClkMux I__11773 (
            .O(N__49928),
            .I(N__49583));
    ClkMux I__11772 (
            .O(N__49927),
            .I(N__49583));
    ClkMux I__11771 (
            .O(N__49926),
            .I(N__49583));
    ClkMux I__11770 (
            .O(N__49925),
            .I(N__49583));
    ClkMux I__11769 (
            .O(N__49924),
            .I(N__49583));
    ClkMux I__11768 (
            .O(N__49923),
            .I(N__49583));
    ClkMux I__11767 (
            .O(N__49922),
            .I(N__49583));
    ClkMux I__11766 (
            .O(N__49921),
            .I(N__49583));
    ClkMux I__11765 (
            .O(N__49920),
            .I(N__49583));
    ClkMux I__11764 (
            .O(N__49919),
            .I(N__49583));
    ClkMux I__11763 (
            .O(N__49918),
            .I(N__49583));
    ClkMux I__11762 (
            .O(N__49917),
            .I(N__49583));
    ClkMux I__11761 (
            .O(N__49916),
            .I(N__49583));
    ClkMux I__11760 (
            .O(N__49915),
            .I(N__49583));
    ClkMux I__11759 (
            .O(N__49914),
            .I(N__49583));
    ClkMux I__11758 (
            .O(N__49913),
            .I(N__49583));
    ClkMux I__11757 (
            .O(N__49912),
            .I(N__49583));
    ClkMux I__11756 (
            .O(N__49911),
            .I(N__49583));
    ClkMux I__11755 (
            .O(N__49910),
            .I(N__49583));
    ClkMux I__11754 (
            .O(N__49909),
            .I(N__49583));
    ClkMux I__11753 (
            .O(N__49908),
            .I(N__49583));
    ClkMux I__11752 (
            .O(N__49907),
            .I(N__49583));
    ClkMux I__11751 (
            .O(N__49906),
            .I(N__49583));
    ClkMux I__11750 (
            .O(N__49905),
            .I(N__49583));
    ClkMux I__11749 (
            .O(N__49904),
            .I(N__49583));
    ClkMux I__11748 (
            .O(N__49903),
            .I(N__49583));
    ClkMux I__11747 (
            .O(N__49902),
            .I(N__49583));
    ClkMux I__11746 (
            .O(N__49901),
            .I(N__49583));
    ClkMux I__11745 (
            .O(N__49900),
            .I(N__49583));
    ClkMux I__11744 (
            .O(N__49899),
            .I(N__49583));
    Glb2LocalMux I__11743 (
            .O(N__49896),
            .I(N__49583));
    ClkMux I__11742 (
            .O(N__49895),
            .I(N__49583));
    ClkMux I__11741 (
            .O(N__49894),
            .I(N__49583));
    GlobalMux I__11740 (
            .O(N__49583),
            .I(clock_output_0));
    InMux I__11739 (
            .O(N__49580),
            .I(N__49570));
    InMux I__11738 (
            .O(N__49579),
            .I(N__49570));
    InMux I__11737 (
            .O(N__49578),
            .I(N__49570));
    CEMux I__11736 (
            .O(N__49577),
            .I(N__49567));
    LocalMux I__11735 (
            .O(N__49570),
            .I(N__49560));
    LocalMux I__11734 (
            .O(N__49567),
            .I(N__49557));
    CEMux I__11733 (
            .O(N__49566),
            .I(N__49554));
    CEMux I__11732 (
            .O(N__49565),
            .I(N__49551));
    CEMux I__11731 (
            .O(N__49564),
            .I(N__49545));
    CEMux I__11730 (
            .O(N__49563),
            .I(N__49539));
    Span4Mux_v I__11729 (
            .O(N__49560),
            .I(N__49530));
    Span4Mux_h I__11728 (
            .O(N__49557),
            .I(N__49530));
    LocalMux I__11727 (
            .O(N__49554),
            .I(N__49530));
    LocalMux I__11726 (
            .O(N__49551),
            .I(N__49530));
    CEMux I__11725 (
            .O(N__49550),
            .I(N__49517));
    CEMux I__11724 (
            .O(N__49549),
            .I(N__49514));
    CEMux I__11723 (
            .O(N__49548),
            .I(N__49511));
    LocalMux I__11722 (
            .O(N__49545),
            .I(N__49508));
    CEMux I__11721 (
            .O(N__49544),
            .I(N__49505));
    CEMux I__11720 (
            .O(N__49543),
            .I(N__49502));
    CEMux I__11719 (
            .O(N__49542),
            .I(N__49497));
    LocalMux I__11718 (
            .O(N__49539),
            .I(N__49494));
    Span4Mux_v I__11717 (
            .O(N__49530),
            .I(N__49491));
    InMux I__11716 (
            .O(N__49529),
            .I(N__49482));
    InMux I__11715 (
            .O(N__49528),
            .I(N__49482));
    InMux I__11714 (
            .O(N__49527),
            .I(N__49482));
    InMux I__11713 (
            .O(N__49526),
            .I(N__49482));
    InMux I__11712 (
            .O(N__49525),
            .I(N__49473));
    InMux I__11711 (
            .O(N__49524),
            .I(N__49473));
    InMux I__11710 (
            .O(N__49523),
            .I(N__49473));
    InMux I__11709 (
            .O(N__49522),
            .I(N__49473));
    CEMux I__11708 (
            .O(N__49521),
            .I(N__49466));
    CEMux I__11707 (
            .O(N__49520),
            .I(N__49457));
    LocalMux I__11706 (
            .O(N__49517),
            .I(N__49454));
    LocalMux I__11705 (
            .O(N__49514),
            .I(N__49451));
    LocalMux I__11704 (
            .O(N__49511),
            .I(N__49448));
    Span4Mux_h I__11703 (
            .O(N__49508),
            .I(N__49443));
    LocalMux I__11702 (
            .O(N__49505),
            .I(N__49443));
    LocalMux I__11701 (
            .O(N__49502),
            .I(N__49440));
    CEMux I__11700 (
            .O(N__49501),
            .I(N__49437));
    CEMux I__11699 (
            .O(N__49500),
            .I(N__49430));
    LocalMux I__11698 (
            .O(N__49497),
            .I(N__49426));
    Span4Mux_h I__11697 (
            .O(N__49494),
            .I(N__49417));
    Span4Mux_h I__11696 (
            .O(N__49491),
            .I(N__49417));
    LocalMux I__11695 (
            .O(N__49482),
            .I(N__49417));
    LocalMux I__11694 (
            .O(N__49473),
            .I(N__49417));
    InMux I__11693 (
            .O(N__49472),
            .I(N__49408));
    InMux I__11692 (
            .O(N__49471),
            .I(N__49408));
    InMux I__11691 (
            .O(N__49470),
            .I(N__49408));
    InMux I__11690 (
            .O(N__49469),
            .I(N__49408));
    LocalMux I__11689 (
            .O(N__49466),
            .I(N__49405));
    CEMux I__11688 (
            .O(N__49465),
            .I(N__49402));
    InMux I__11687 (
            .O(N__49464),
            .I(N__49393));
    InMux I__11686 (
            .O(N__49463),
            .I(N__49393));
    InMux I__11685 (
            .O(N__49462),
            .I(N__49393));
    InMux I__11684 (
            .O(N__49461),
            .I(N__49393));
    CEMux I__11683 (
            .O(N__49460),
            .I(N__49390));
    LocalMux I__11682 (
            .O(N__49457),
            .I(N__49378));
    Span4Mux_h I__11681 (
            .O(N__49454),
            .I(N__49378));
    Span4Mux_h I__11680 (
            .O(N__49451),
            .I(N__49378));
    Span4Mux_h I__11679 (
            .O(N__49448),
            .I(N__49378));
    Span4Mux_v I__11678 (
            .O(N__49443),
            .I(N__49375));
    Span4Mux_v I__11677 (
            .O(N__49440),
            .I(N__49372));
    LocalMux I__11676 (
            .O(N__49437),
            .I(N__49369));
    InMux I__11675 (
            .O(N__49436),
            .I(N__49360));
    InMux I__11674 (
            .O(N__49435),
            .I(N__49360));
    InMux I__11673 (
            .O(N__49434),
            .I(N__49360));
    InMux I__11672 (
            .O(N__49433),
            .I(N__49360));
    LocalMux I__11671 (
            .O(N__49430),
            .I(N__49353));
    InMux I__11670 (
            .O(N__49429),
            .I(N__49350));
    Span4Mux_v I__11669 (
            .O(N__49426),
            .I(N__49347));
    Span4Mux_v I__11668 (
            .O(N__49417),
            .I(N__49342));
    LocalMux I__11667 (
            .O(N__49408),
            .I(N__49342));
    Span4Mux_s2_v I__11666 (
            .O(N__49405),
            .I(N__49339));
    LocalMux I__11665 (
            .O(N__49402),
            .I(N__49334));
    LocalMux I__11664 (
            .O(N__49393),
            .I(N__49334));
    LocalMux I__11663 (
            .O(N__49390),
            .I(N__49331));
    InMux I__11662 (
            .O(N__49389),
            .I(N__49324));
    InMux I__11661 (
            .O(N__49388),
            .I(N__49324));
    InMux I__11660 (
            .O(N__49387),
            .I(N__49324));
    Span4Mux_v I__11659 (
            .O(N__49378),
            .I(N__49321));
    Span4Mux_s1_v I__11658 (
            .O(N__49375),
            .I(N__49316));
    Span4Mux_h I__11657 (
            .O(N__49372),
            .I(N__49316));
    Span4Mux_h I__11656 (
            .O(N__49369),
            .I(N__49311));
    LocalMux I__11655 (
            .O(N__49360),
            .I(N__49311));
    InMux I__11654 (
            .O(N__49359),
            .I(N__49302));
    InMux I__11653 (
            .O(N__49358),
            .I(N__49302));
    InMux I__11652 (
            .O(N__49357),
            .I(N__49302));
    InMux I__11651 (
            .O(N__49356),
            .I(N__49302));
    Span4Mux_v I__11650 (
            .O(N__49353),
            .I(N__49297));
    LocalMux I__11649 (
            .O(N__49350),
            .I(N__49297));
    Span4Mux_h I__11648 (
            .O(N__49347),
            .I(N__49288));
    Span4Mux_v I__11647 (
            .O(N__49342),
            .I(N__49288));
    Span4Mux_h I__11646 (
            .O(N__49339),
            .I(N__49288));
    Span4Mux_h I__11645 (
            .O(N__49334),
            .I(N__49288));
    Odrv12 I__11644 (
            .O(N__49331),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__11643 (
            .O(N__49324),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11642 (
            .O(N__49321),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11641 (
            .O(N__49316),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11640 (
            .O(N__49311),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__11639 (
            .O(N__49302),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11638 (
            .O(N__49297),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11637 (
            .O(N__49288),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__11636 (
            .O(N__49271),
            .I(N__49265));
    InMux I__11635 (
            .O(N__49270),
            .I(N__49262));
    InMux I__11634 (
            .O(N__49269),
            .I(N__49259));
    InMux I__11633 (
            .O(N__49268),
            .I(N__49256));
    LocalMux I__11632 (
            .O(N__49265),
            .I(N__49253));
    LocalMux I__11631 (
            .O(N__49262),
            .I(N__49250));
    LocalMux I__11630 (
            .O(N__49259),
            .I(N__49247));
    LocalMux I__11629 (
            .O(N__49256),
            .I(N__49241));
    Glb2LocalMux I__11628 (
            .O(N__49253),
            .I(N__48767));
    Glb2LocalMux I__11627 (
            .O(N__49250),
            .I(N__48767));
    Glb2LocalMux I__11626 (
            .O(N__49247),
            .I(N__48767));
    SRMux I__11625 (
            .O(N__49246),
            .I(N__48767));
    SRMux I__11624 (
            .O(N__49245),
            .I(N__48767));
    SRMux I__11623 (
            .O(N__49244),
            .I(N__48767));
    Glb2LocalMux I__11622 (
            .O(N__49241),
            .I(N__48767));
    SRMux I__11621 (
            .O(N__49240),
            .I(N__48767));
    SRMux I__11620 (
            .O(N__49239),
            .I(N__48767));
    SRMux I__11619 (
            .O(N__49238),
            .I(N__48767));
    SRMux I__11618 (
            .O(N__49237),
            .I(N__48767));
    SRMux I__11617 (
            .O(N__49236),
            .I(N__48767));
    SRMux I__11616 (
            .O(N__49235),
            .I(N__48767));
    SRMux I__11615 (
            .O(N__49234),
            .I(N__48767));
    SRMux I__11614 (
            .O(N__49233),
            .I(N__48767));
    SRMux I__11613 (
            .O(N__49232),
            .I(N__48767));
    SRMux I__11612 (
            .O(N__49231),
            .I(N__48767));
    SRMux I__11611 (
            .O(N__49230),
            .I(N__48767));
    SRMux I__11610 (
            .O(N__49229),
            .I(N__48767));
    SRMux I__11609 (
            .O(N__49228),
            .I(N__48767));
    SRMux I__11608 (
            .O(N__49227),
            .I(N__48767));
    SRMux I__11607 (
            .O(N__49226),
            .I(N__48767));
    SRMux I__11606 (
            .O(N__49225),
            .I(N__48767));
    SRMux I__11605 (
            .O(N__49224),
            .I(N__48767));
    SRMux I__11604 (
            .O(N__49223),
            .I(N__48767));
    SRMux I__11603 (
            .O(N__49222),
            .I(N__48767));
    SRMux I__11602 (
            .O(N__49221),
            .I(N__48767));
    SRMux I__11601 (
            .O(N__49220),
            .I(N__48767));
    SRMux I__11600 (
            .O(N__49219),
            .I(N__48767));
    SRMux I__11599 (
            .O(N__49218),
            .I(N__48767));
    SRMux I__11598 (
            .O(N__49217),
            .I(N__48767));
    SRMux I__11597 (
            .O(N__49216),
            .I(N__48767));
    SRMux I__11596 (
            .O(N__49215),
            .I(N__48767));
    SRMux I__11595 (
            .O(N__49214),
            .I(N__48767));
    SRMux I__11594 (
            .O(N__49213),
            .I(N__48767));
    SRMux I__11593 (
            .O(N__49212),
            .I(N__48767));
    SRMux I__11592 (
            .O(N__49211),
            .I(N__48767));
    SRMux I__11591 (
            .O(N__49210),
            .I(N__48767));
    SRMux I__11590 (
            .O(N__49209),
            .I(N__48767));
    SRMux I__11589 (
            .O(N__49208),
            .I(N__48767));
    SRMux I__11588 (
            .O(N__49207),
            .I(N__48767));
    SRMux I__11587 (
            .O(N__49206),
            .I(N__48767));
    SRMux I__11586 (
            .O(N__49205),
            .I(N__48767));
    SRMux I__11585 (
            .O(N__49204),
            .I(N__48767));
    SRMux I__11584 (
            .O(N__49203),
            .I(N__48767));
    SRMux I__11583 (
            .O(N__49202),
            .I(N__48767));
    SRMux I__11582 (
            .O(N__49201),
            .I(N__48767));
    SRMux I__11581 (
            .O(N__49200),
            .I(N__48767));
    SRMux I__11580 (
            .O(N__49199),
            .I(N__48767));
    SRMux I__11579 (
            .O(N__49198),
            .I(N__48767));
    SRMux I__11578 (
            .O(N__49197),
            .I(N__48767));
    SRMux I__11577 (
            .O(N__49196),
            .I(N__48767));
    SRMux I__11576 (
            .O(N__49195),
            .I(N__48767));
    SRMux I__11575 (
            .O(N__49194),
            .I(N__48767));
    SRMux I__11574 (
            .O(N__49193),
            .I(N__48767));
    SRMux I__11573 (
            .O(N__49192),
            .I(N__48767));
    SRMux I__11572 (
            .O(N__49191),
            .I(N__48767));
    SRMux I__11571 (
            .O(N__49190),
            .I(N__48767));
    SRMux I__11570 (
            .O(N__49189),
            .I(N__48767));
    SRMux I__11569 (
            .O(N__49188),
            .I(N__48767));
    SRMux I__11568 (
            .O(N__49187),
            .I(N__48767));
    SRMux I__11567 (
            .O(N__49186),
            .I(N__48767));
    SRMux I__11566 (
            .O(N__49185),
            .I(N__48767));
    SRMux I__11565 (
            .O(N__49184),
            .I(N__48767));
    SRMux I__11564 (
            .O(N__49183),
            .I(N__48767));
    SRMux I__11563 (
            .O(N__49182),
            .I(N__48767));
    SRMux I__11562 (
            .O(N__49181),
            .I(N__48767));
    SRMux I__11561 (
            .O(N__49180),
            .I(N__48767));
    SRMux I__11560 (
            .O(N__49179),
            .I(N__48767));
    SRMux I__11559 (
            .O(N__49178),
            .I(N__48767));
    SRMux I__11558 (
            .O(N__49177),
            .I(N__48767));
    SRMux I__11557 (
            .O(N__49176),
            .I(N__48767));
    SRMux I__11556 (
            .O(N__49175),
            .I(N__48767));
    SRMux I__11555 (
            .O(N__49174),
            .I(N__48767));
    SRMux I__11554 (
            .O(N__49173),
            .I(N__48767));
    SRMux I__11553 (
            .O(N__49172),
            .I(N__48767));
    SRMux I__11552 (
            .O(N__49171),
            .I(N__48767));
    SRMux I__11551 (
            .O(N__49170),
            .I(N__48767));
    SRMux I__11550 (
            .O(N__49169),
            .I(N__48767));
    SRMux I__11549 (
            .O(N__49168),
            .I(N__48767));
    SRMux I__11548 (
            .O(N__49167),
            .I(N__48767));
    SRMux I__11547 (
            .O(N__49166),
            .I(N__48767));
    SRMux I__11546 (
            .O(N__49165),
            .I(N__48767));
    SRMux I__11545 (
            .O(N__49164),
            .I(N__48767));
    SRMux I__11544 (
            .O(N__49163),
            .I(N__48767));
    SRMux I__11543 (
            .O(N__49162),
            .I(N__48767));
    SRMux I__11542 (
            .O(N__49161),
            .I(N__48767));
    SRMux I__11541 (
            .O(N__49160),
            .I(N__48767));
    SRMux I__11540 (
            .O(N__49159),
            .I(N__48767));
    SRMux I__11539 (
            .O(N__49158),
            .I(N__48767));
    SRMux I__11538 (
            .O(N__49157),
            .I(N__48767));
    SRMux I__11537 (
            .O(N__49156),
            .I(N__48767));
    SRMux I__11536 (
            .O(N__49155),
            .I(N__48767));
    SRMux I__11535 (
            .O(N__49154),
            .I(N__48767));
    SRMux I__11534 (
            .O(N__49153),
            .I(N__48767));
    SRMux I__11533 (
            .O(N__49152),
            .I(N__48767));
    SRMux I__11532 (
            .O(N__49151),
            .I(N__48767));
    SRMux I__11531 (
            .O(N__49150),
            .I(N__48767));
    SRMux I__11530 (
            .O(N__49149),
            .I(N__48767));
    SRMux I__11529 (
            .O(N__49148),
            .I(N__48767));
    SRMux I__11528 (
            .O(N__49147),
            .I(N__48767));
    SRMux I__11527 (
            .O(N__49146),
            .I(N__48767));
    SRMux I__11526 (
            .O(N__49145),
            .I(N__48767));
    SRMux I__11525 (
            .O(N__49144),
            .I(N__48767));
    SRMux I__11524 (
            .O(N__49143),
            .I(N__48767));
    SRMux I__11523 (
            .O(N__49142),
            .I(N__48767));
    SRMux I__11522 (
            .O(N__49141),
            .I(N__48767));
    SRMux I__11521 (
            .O(N__49140),
            .I(N__48767));
    SRMux I__11520 (
            .O(N__49139),
            .I(N__48767));
    SRMux I__11519 (
            .O(N__49138),
            .I(N__48767));
    SRMux I__11518 (
            .O(N__49137),
            .I(N__48767));
    SRMux I__11517 (
            .O(N__49136),
            .I(N__48767));
    SRMux I__11516 (
            .O(N__49135),
            .I(N__48767));
    SRMux I__11515 (
            .O(N__49134),
            .I(N__48767));
    SRMux I__11514 (
            .O(N__49133),
            .I(N__48767));
    SRMux I__11513 (
            .O(N__49132),
            .I(N__48767));
    SRMux I__11512 (
            .O(N__49131),
            .I(N__48767));
    SRMux I__11511 (
            .O(N__49130),
            .I(N__48767));
    SRMux I__11510 (
            .O(N__49129),
            .I(N__48767));
    SRMux I__11509 (
            .O(N__49128),
            .I(N__48767));
    SRMux I__11508 (
            .O(N__49127),
            .I(N__48767));
    SRMux I__11507 (
            .O(N__49126),
            .I(N__48767));
    SRMux I__11506 (
            .O(N__49125),
            .I(N__48767));
    SRMux I__11505 (
            .O(N__49124),
            .I(N__48767));
    SRMux I__11504 (
            .O(N__49123),
            .I(N__48767));
    SRMux I__11503 (
            .O(N__49122),
            .I(N__48767));
    SRMux I__11502 (
            .O(N__49121),
            .I(N__48767));
    SRMux I__11501 (
            .O(N__49120),
            .I(N__48767));
    SRMux I__11500 (
            .O(N__49119),
            .I(N__48767));
    SRMux I__11499 (
            .O(N__49118),
            .I(N__48767));
    SRMux I__11498 (
            .O(N__49117),
            .I(N__48767));
    SRMux I__11497 (
            .O(N__49116),
            .I(N__48767));
    SRMux I__11496 (
            .O(N__49115),
            .I(N__48767));
    SRMux I__11495 (
            .O(N__49114),
            .I(N__48767));
    SRMux I__11494 (
            .O(N__49113),
            .I(N__48767));
    SRMux I__11493 (
            .O(N__49112),
            .I(N__48767));
    SRMux I__11492 (
            .O(N__49111),
            .I(N__48767));
    SRMux I__11491 (
            .O(N__49110),
            .I(N__48767));
    SRMux I__11490 (
            .O(N__49109),
            .I(N__48767));
    SRMux I__11489 (
            .O(N__49108),
            .I(N__48767));
    SRMux I__11488 (
            .O(N__49107),
            .I(N__48767));
    SRMux I__11487 (
            .O(N__49106),
            .I(N__48767));
    SRMux I__11486 (
            .O(N__49105),
            .I(N__48767));
    SRMux I__11485 (
            .O(N__49104),
            .I(N__48767));
    SRMux I__11484 (
            .O(N__49103),
            .I(N__48767));
    SRMux I__11483 (
            .O(N__49102),
            .I(N__48767));
    SRMux I__11482 (
            .O(N__49101),
            .I(N__48767));
    SRMux I__11481 (
            .O(N__49100),
            .I(N__48767));
    SRMux I__11480 (
            .O(N__49099),
            .I(N__48767));
    SRMux I__11479 (
            .O(N__49098),
            .I(N__48767));
    SRMux I__11478 (
            .O(N__49097),
            .I(N__48767));
    SRMux I__11477 (
            .O(N__49096),
            .I(N__48767));
    SRMux I__11476 (
            .O(N__49095),
            .I(N__48767));
    SRMux I__11475 (
            .O(N__49094),
            .I(N__48767));
    SRMux I__11474 (
            .O(N__49093),
            .I(N__48767));
    SRMux I__11473 (
            .O(N__49092),
            .I(N__48767));
    SRMux I__11472 (
            .O(N__49091),
            .I(N__48767));
    SRMux I__11471 (
            .O(N__49090),
            .I(N__48767));
    SRMux I__11470 (
            .O(N__49089),
            .I(N__48767));
    SRMux I__11469 (
            .O(N__49088),
            .I(N__48767));
    GlobalMux I__11468 (
            .O(N__48767),
            .I(N__48764));
    gio2CtrlBuf I__11467 (
            .O(N__48764),
            .I(red_c_g));
    InMux I__11466 (
            .O(N__48761),
            .I(N__48754));
    InMux I__11465 (
            .O(N__48760),
            .I(N__48754));
    InMux I__11464 (
            .O(N__48759),
            .I(N__48751));
    LocalMux I__11463 (
            .O(N__48754),
            .I(N__48748));
    LocalMux I__11462 (
            .O(N__48751),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv12 I__11461 (
            .O(N__48748),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__11460 (
            .O(N__48743),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__11459 (
            .O(N__48740),
            .I(N__48736));
    CascadeMux I__11458 (
            .O(N__48739),
            .I(N__48733));
    InMux I__11457 (
            .O(N__48736),
            .I(N__48727));
    InMux I__11456 (
            .O(N__48733),
            .I(N__48727));
    InMux I__11455 (
            .O(N__48732),
            .I(N__48724));
    LocalMux I__11454 (
            .O(N__48727),
            .I(N__48721));
    LocalMux I__11453 (
            .O(N__48724),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv12 I__11452 (
            .O(N__48721),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__11451 (
            .O(N__48716),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__11450 (
            .O(N__48713),
            .I(N__48709));
    InMux I__11449 (
            .O(N__48712),
            .I(N__48705));
    InMux I__11448 (
            .O(N__48709),
            .I(N__48702));
    InMux I__11447 (
            .O(N__48708),
            .I(N__48699));
    LocalMux I__11446 (
            .O(N__48705),
            .I(N__48694));
    LocalMux I__11445 (
            .O(N__48702),
            .I(N__48694));
    LocalMux I__11444 (
            .O(N__48699),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv12 I__11443 (
            .O(N__48694),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__11442 (
            .O(N__48689),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__11441 (
            .O(N__48686),
            .I(N__48683));
    InMux I__11440 (
            .O(N__48683),
            .I(N__48678));
    InMux I__11439 (
            .O(N__48682),
            .I(N__48675));
    InMux I__11438 (
            .O(N__48681),
            .I(N__48672));
    LocalMux I__11437 (
            .O(N__48678),
            .I(N__48667));
    LocalMux I__11436 (
            .O(N__48675),
            .I(N__48667));
    LocalMux I__11435 (
            .O(N__48672),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv12 I__11434 (
            .O(N__48667),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__11433 (
            .O(N__48662),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__11432 (
            .O(N__48659),
            .I(N__48655));
    CascadeMux I__11431 (
            .O(N__48658),
            .I(N__48652));
    InMux I__11430 (
            .O(N__48655),
            .I(N__48647));
    InMux I__11429 (
            .O(N__48652),
            .I(N__48647));
    LocalMux I__11428 (
            .O(N__48647),
            .I(N__48643));
    InMux I__11427 (
            .O(N__48646),
            .I(N__48640));
    Span4Mux_v I__11426 (
            .O(N__48643),
            .I(N__48637));
    LocalMux I__11425 (
            .O(N__48640),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__11424 (
            .O(N__48637),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__11423 (
            .O(N__48632),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__11422 (
            .O(N__48629),
            .I(N__48622));
    InMux I__11421 (
            .O(N__48628),
            .I(N__48622));
    InMux I__11420 (
            .O(N__48627),
            .I(N__48619));
    LocalMux I__11419 (
            .O(N__48622),
            .I(N__48616));
    LocalMux I__11418 (
            .O(N__48619),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv12 I__11417 (
            .O(N__48616),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__11416 (
            .O(N__48611),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__11415 (
            .O(N__48608),
            .I(N__48605));
    InMux I__11414 (
            .O(N__48605),
            .I(N__48601));
    InMux I__11413 (
            .O(N__48604),
            .I(N__48598));
    LocalMux I__11412 (
            .O(N__48601),
            .I(N__48592));
    LocalMux I__11411 (
            .O(N__48598),
            .I(N__48592));
    InMux I__11410 (
            .O(N__48597),
            .I(N__48589));
    Span4Mux_v I__11409 (
            .O(N__48592),
            .I(N__48586));
    LocalMux I__11408 (
            .O(N__48589),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__11407 (
            .O(N__48586),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__11406 (
            .O(N__48581),
            .I(bfn_18_26_0_));
    CascadeMux I__11405 (
            .O(N__48578),
            .I(N__48574));
    InMux I__11404 (
            .O(N__48577),
            .I(N__48571));
    InMux I__11403 (
            .O(N__48574),
            .I(N__48568));
    LocalMux I__11402 (
            .O(N__48571),
            .I(N__48562));
    LocalMux I__11401 (
            .O(N__48568),
            .I(N__48562));
    InMux I__11400 (
            .O(N__48567),
            .I(N__48559));
    Span4Mux_v I__11399 (
            .O(N__48562),
            .I(N__48556));
    LocalMux I__11398 (
            .O(N__48559),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__11397 (
            .O(N__48556),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__11396 (
            .O(N__48551),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__11395 (
            .O(N__48548),
            .I(N__48545));
    InMux I__11394 (
            .O(N__48545),
            .I(N__48541));
    InMux I__11393 (
            .O(N__48544),
            .I(N__48538));
    LocalMux I__11392 (
            .O(N__48541),
            .I(N__48532));
    LocalMux I__11391 (
            .O(N__48538),
            .I(N__48532));
    InMux I__11390 (
            .O(N__48537),
            .I(N__48529));
    Span4Mux_v I__11389 (
            .O(N__48532),
            .I(N__48526));
    LocalMux I__11388 (
            .O(N__48529),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__11387 (
            .O(N__48526),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__11386 (
            .O(N__48521),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__11385 (
            .O(N__48518),
            .I(N__48512));
    InMux I__11384 (
            .O(N__48517),
            .I(N__48512));
    LocalMux I__11383 (
            .O(N__48512),
            .I(N__48508));
    InMux I__11382 (
            .O(N__48511),
            .I(N__48505));
    Span4Mux_h I__11381 (
            .O(N__48508),
            .I(N__48502));
    LocalMux I__11380 (
            .O(N__48505),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__11379 (
            .O(N__48502),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__11378 (
            .O(N__48497),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__11377 (
            .O(N__48494),
            .I(N__48488));
    InMux I__11376 (
            .O(N__48493),
            .I(N__48488));
    LocalMux I__11375 (
            .O(N__48488),
            .I(N__48484));
    InMux I__11374 (
            .O(N__48487),
            .I(N__48481));
    Span4Mux_h I__11373 (
            .O(N__48484),
            .I(N__48478));
    LocalMux I__11372 (
            .O(N__48481),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__11371 (
            .O(N__48478),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__11370 (
            .O(N__48473),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__11369 (
            .O(N__48470),
            .I(N__48466));
    CascadeMux I__11368 (
            .O(N__48469),
            .I(N__48463));
    InMux I__11367 (
            .O(N__48466),
            .I(N__48458));
    InMux I__11366 (
            .O(N__48463),
            .I(N__48458));
    LocalMux I__11365 (
            .O(N__48458),
            .I(N__48454));
    InMux I__11364 (
            .O(N__48457),
            .I(N__48451));
    Span4Mux_v I__11363 (
            .O(N__48454),
            .I(N__48448));
    LocalMux I__11362 (
            .O(N__48451),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__11361 (
            .O(N__48448),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__11360 (
            .O(N__48443),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__11359 (
            .O(N__48440),
            .I(N__48436));
    CascadeMux I__11358 (
            .O(N__48439),
            .I(N__48433));
    InMux I__11357 (
            .O(N__48436),
            .I(N__48428));
    InMux I__11356 (
            .O(N__48433),
            .I(N__48428));
    LocalMux I__11355 (
            .O(N__48428),
            .I(N__48424));
    InMux I__11354 (
            .O(N__48427),
            .I(N__48421));
    Span4Mux_h I__11353 (
            .O(N__48424),
            .I(N__48418));
    LocalMux I__11352 (
            .O(N__48421),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__11351 (
            .O(N__48418),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__11350 (
            .O(N__48413),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__11349 (
            .O(N__48410),
            .I(N__48404));
    InMux I__11348 (
            .O(N__48409),
            .I(N__48404));
    LocalMux I__11347 (
            .O(N__48404),
            .I(N__48400));
    InMux I__11346 (
            .O(N__48403),
            .I(N__48397));
    Span4Mux_v I__11345 (
            .O(N__48400),
            .I(N__48394));
    LocalMux I__11344 (
            .O(N__48397),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__11343 (
            .O(N__48394),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__11342 (
            .O(N__48389),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    CascadeMux I__11341 (
            .O(N__48386),
            .I(N__48383));
    InMux I__11340 (
            .O(N__48383),
            .I(N__48379));
    InMux I__11339 (
            .O(N__48382),
            .I(N__48376));
    LocalMux I__11338 (
            .O(N__48379),
            .I(N__48370));
    LocalMux I__11337 (
            .O(N__48376),
            .I(N__48370));
    InMux I__11336 (
            .O(N__48375),
            .I(N__48367));
    Span4Mux_v I__11335 (
            .O(N__48370),
            .I(N__48364));
    LocalMux I__11334 (
            .O(N__48367),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__11333 (
            .O(N__48364),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__11332 (
            .O(N__48359),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__11331 (
            .O(N__48356),
            .I(N__48352));
    CascadeMux I__11330 (
            .O(N__48355),
            .I(N__48349));
    InMux I__11329 (
            .O(N__48352),
            .I(N__48346));
    InMux I__11328 (
            .O(N__48349),
            .I(N__48343));
    LocalMux I__11327 (
            .O(N__48346),
            .I(N__48337));
    LocalMux I__11326 (
            .O(N__48343),
            .I(N__48337));
    InMux I__11325 (
            .O(N__48342),
            .I(N__48334));
    Span4Mux_v I__11324 (
            .O(N__48337),
            .I(N__48331));
    LocalMux I__11323 (
            .O(N__48334),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__11322 (
            .O(N__48331),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__11321 (
            .O(N__48326),
            .I(bfn_18_25_0_));
    InMux I__11320 (
            .O(N__48323),
            .I(N__48319));
    InMux I__11319 (
            .O(N__48322),
            .I(N__48316));
    LocalMux I__11318 (
            .O(N__48319),
            .I(N__48310));
    LocalMux I__11317 (
            .O(N__48316),
            .I(N__48310));
    InMux I__11316 (
            .O(N__48315),
            .I(N__48307));
    Span4Mux_v I__11315 (
            .O(N__48310),
            .I(N__48304));
    LocalMux I__11314 (
            .O(N__48307),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__11313 (
            .O(N__48304),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__11312 (
            .O(N__48299),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__11311 (
            .O(N__48296),
            .I(N__48293));
    LocalMux I__11310 (
            .O(N__48293),
            .I(N__48289));
    CascadeMux I__11309 (
            .O(N__48292),
            .I(N__48286));
    Span4Mux_v I__11308 (
            .O(N__48289),
            .I(N__48283));
    InMux I__11307 (
            .O(N__48286),
            .I(N__48280));
    Span4Mux_v I__11306 (
            .O(N__48283),
            .I(N__48277));
    LocalMux I__11305 (
            .O(N__48280),
            .I(N__48273));
    Span4Mux_v I__11304 (
            .O(N__48277),
            .I(N__48270));
    InMux I__11303 (
            .O(N__48276),
            .I(N__48267));
    Span4Mux_h I__11302 (
            .O(N__48273),
            .I(N__48264));
    Odrv4 I__11301 (
            .O(N__48270),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__11300 (
            .O(N__48267),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__11299 (
            .O(N__48264),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__11298 (
            .O(N__48257),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__11297 (
            .O(N__48254),
            .I(N__48247));
    InMux I__11296 (
            .O(N__48253),
            .I(N__48247));
    InMux I__11295 (
            .O(N__48252),
            .I(N__48244));
    LocalMux I__11294 (
            .O(N__48247),
            .I(N__48241));
    LocalMux I__11293 (
            .O(N__48244),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__11292 (
            .O(N__48241),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__11291 (
            .O(N__48236),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__11290 (
            .O(N__48233),
            .I(N__48226));
    InMux I__11289 (
            .O(N__48232),
            .I(N__48226));
    InMux I__11288 (
            .O(N__48231),
            .I(N__48223));
    LocalMux I__11287 (
            .O(N__48226),
            .I(N__48220));
    LocalMux I__11286 (
            .O(N__48223),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv12 I__11285 (
            .O(N__48220),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__11284 (
            .O(N__48215),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__11283 (
            .O(N__48212),
            .I(N__48208));
    InMux I__11282 (
            .O(N__48211),
            .I(N__48205));
    InMux I__11281 (
            .O(N__48208),
            .I(N__48202));
    LocalMux I__11280 (
            .O(N__48205),
            .I(N__48196));
    LocalMux I__11279 (
            .O(N__48202),
            .I(N__48196));
    InMux I__11278 (
            .O(N__48201),
            .I(N__48193));
    Span4Mux_h I__11277 (
            .O(N__48196),
            .I(N__48190));
    LocalMux I__11276 (
            .O(N__48193),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__11275 (
            .O(N__48190),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__11274 (
            .O(N__48185),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__11273 (
            .O(N__48182),
            .I(N__48178));
    InMux I__11272 (
            .O(N__48181),
            .I(N__48175));
    InMux I__11271 (
            .O(N__48178),
            .I(N__48172));
    LocalMux I__11270 (
            .O(N__48175),
            .I(N__48166));
    LocalMux I__11269 (
            .O(N__48172),
            .I(N__48166));
    InMux I__11268 (
            .O(N__48171),
            .I(N__48163));
    Span4Mux_h I__11267 (
            .O(N__48166),
            .I(N__48160));
    LocalMux I__11266 (
            .O(N__48163),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__11265 (
            .O(N__48160),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__11264 (
            .O(N__48155),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__11263 (
            .O(N__48152),
            .I(N__48148));
    CascadeMux I__11262 (
            .O(N__48151),
            .I(N__48145));
    InMux I__11261 (
            .O(N__48148),
            .I(N__48140));
    InMux I__11260 (
            .O(N__48145),
            .I(N__48140));
    LocalMux I__11259 (
            .O(N__48140),
            .I(N__48136));
    InMux I__11258 (
            .O(N__48139),
            .I(N__48133));
    Span4Mux_v I__11257 (
            .O(N__48136),
            .I(N__48130));
    LocalMux I__11256 (
            .O(N__48133),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__11255 (
            .O(N__48130),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__11254 (
            .O(N__48125),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    CascadeMux I__11253 (
            .O(N__48122),
            .I(N__48118));
    CascadeMux I__11252 (
            .O(N__48121),
            .I(N__48115));
    InMux I__11251 (
            .O(N__48118),
            .I(N__48110));
    InMux I__11250 (
            .O(N__48115),
            .I(N__48110));
    LocalMux I__11249 (
            .O(N__48110),
            .I(N__48106));
    InMux I__11248 (
            .O(N__48109),
            .I(N__48103));
    Span4Mux_v I__11247 (
            .O(N__48106),
            .I(N__48100));
    LocalMux I__11246 (
            .O(N__48103),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__11245 (
            .O(N__48100),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__11244 (
            .O(N__48095),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__11243 (
            .O(N__48092),
            .I(N__48089));
    InMux I__11242 (
            .O(N__48089),
            .I(N__48085));
    InMux I__11241 (
            .O(N__48088),
            .I(N__48082));
    LocalMux I__11240 (
            .O(N__48085),
            .I(N__48076));
    LocalMux I__11239 (
            .O(N__48082),
            .I(N__48076));
    InMux I__11238 (
            .O(N__48081),
            .I(N__48073));
    Span4Mux_v I__11237 (
            .O(N__48076),
            .I(N__48070));
    LocalMux I__11236 (
            .O(N__48073),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__11235 (
            .O(N__48070),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__11234 (
            .O(N__48065),
            .I(bfn_18_24_0_));
    InMux I__11233 (
            .O(N__48062),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__11232 (
            .O(N__48059),
            .I(N__48056));
    InMux I__11231 (
            .O(N__48056),
            .I(N__48052));
    CascadeMux I__11230 (
            .O(N__48055),
            .I(N__48049));
    LocalMux I__11229 (
            .O(N__48052),
            .I(N__48046));
    InMux I__11228 (
            .O(N__48049),
            .I(N__48043));
    Span4Mux_h I__11227 (
            .O(N__48046),
            .I(N__48037));
    LocalMux I__11226 (
            .O(N__48043),
            .I(N__48037));
    InMux I__11225 (
            .O(N__48042),
            .I(N__48034));
    Span4Mux_h I__11224 (
            .O(N__48037),
            .I(N__48030));
    LocalMux I__11223 (
            .O(N__48034),
            .I(N__48027));
    InMux I__11222 (
            .O(N__48033),
            .I(N__48024));
    Odrv4 I__11221 (
            .O(N__48030),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__11220 (
            .O(N__48027),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__11219 (
            .O(N__48024),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__11218 (
            .O(N__48017),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__11217 (
            .O(N__48014),
            .I(N__48011));
    InMux I__11216 (
            .O(N__48011),
            .I(N__48007));
    InMux I__11215 (
            .O(N__48010),
            .I(N__48004));
    LocalMux I__11214 (
            .O(N__48007),
            .I(N__48000));
    LocalMux I__11213 (
            .O(N__48004),
            .I(N__47997));
    InMux I__11212 (
            .O(N__48003),
            .I(N__47994));
    Span4Mux_h I__11211 (
            .O(N__48000),
            .I(N__47990));
    Span4Mux_h I__11210 (
            .O(N__47997),
            .I(N__47987));
    LocalMux I__11209 (
            .O(N__47994),
            .I(N__47984));
    InMux I__11208 (
            .O(N__47993),
            .I(N__47981));
    Odrv4 I__11207 (
            .O(N__47990),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__11206 (
            .O(N__47987),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__11205 (
            .O(N__47984),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__11204 (
            .O(N__47981),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__11203 (
            .O(N__47972),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__11202 (
            .O(N__47969),
            .I(N__47965));
    InMux I__11201 (
            .O(N__47968),
            .I(N__47962));
    InMux I__11200 (
            .O(N__47965),
            .I(N__47959));
    LocalMux I__11199 (
            .O(N__47962),
            .I(N__47956));
    LocalMux I__11198 (
            .O(N__47959),
            .I(N__47952));
    Span4Mux_h I__11197 (
            .O(N__47956),
            .I(N__47949));
    InMux I__11196 (
            .O(N__47955),
            .I(N__47946));
    Span4Mux_h I__11195 (
            .O(N__47952),
            .I(N__47942));
    Span4Mux_v I__11194 (
            .O(N__47949),
            .I(N__47937));
    LocalMux I__11193 (
            .O(N__47946),
            .I(N__47937));
    InMux I__11192 (
            .O(N__47945),
            .I(N__47934));
    Odrv4 I__11191 (
            .O(N__47942),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__11190 (
            .O(N__47937),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__11189 (
            .O(N__47934),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__11188 (
            .O(N__47927),
            .I(bfn_18_22_0_));
    CascadeMux I__11187 (
            .O(N__47924),
            .I(N__47920));
    CascadeMux I__11186 (
            .O(N__47923),
            .I(N__47917));
    InMux I__11185 (
            .O(N__47920),
            .I(N__47914));
    InMux I__11184 (
            .O(N__47917),
            .I(N__47911));
    LocalMux I__11183 (
            .O(N__47914),
            .I(N__47907));
    LocalMux I__11182 (
            .O(N__47911),
            .I(N__47904));
    InMux I__11181 (
            .O(N__47910),
            .I(N__47901));
    Span4Mux_h I__11180 (
            .O(N__47907),
            .I(N__47897));
    Span4Mux_h I__11179 (
            .O(N__47904),
            .I(N__47894));
    LocalMux I__11178 (
            .O(N__47901),
            .I(N__47891));
    InMux I__11177 (
            .O(N__47900),
            .I(N__47888));
    Odrv4 I__11176 (
            .O(N__47897),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__11175 (
            .O(N__47894),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__11174 (
            .O(N__47891),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__11173 (
            .O(N__47888),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__11172 (
            .O(N__47879),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__11171 (
            .O(N__47876),
            .I(N__47872));
    InMux I__11170 (
            .O(N__47875),
            .I(N__47869));
    LocalMux I__11169 (
            .O(N__47872),
            .I(N__47863));
    LocalMux I__11168 (
            .O(N__47869),
            .I(N__47863));
    InMux I__11167 (
            .O(N__47868),
            .I(N__47860));
    Span4Mux_v I__11166 (
            .O(N__47863),
            .I(N__47856));
    LocalMux I__11165 (
            .O(N__47860),
            .I(N__47853));
    InMux I__11164 (
            .O(N__47859),
            .I(N__47850));
    Odrv4 I__11163 (
            .O(N__47856),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__11162 (
            .O(N__47853),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__11161 (
            .O(N__47850),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__11160 (
            .O(N__47843),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__11159 (
            .O(N__47840),
            .I(N__47837));
    InMux I__11158 (
            .O(N__47837),
            .I(N__47833));
    CascadeMux I__11157 (
            .O(N__47836),
            .I(N__47830));
    LocalMux I__11156 (
            .O(N__47833),
            .I(N__47827));
    InMux I__11155 (
            .O(N__47830),
            .I(N__47824));
    Span4Mux_v I__11154 (
            .O(N__47827),
            .I(N__47818));
    LocalMux I__11153 (
            .O(N__47824),
            .I(N__47818));
    InMux I__11152 (
            .O(N__47823),
            .I(N__47815));
    Span4Mux_h I__11151 (
            .O(N__47818),
            .I(N__47811));
    LocalMux I__11150 (
            .O(N__47815),
            .I(N__47808));
    InMux I__11149 (
            .O(N__47814),
            .I(N__47805));
    Odrv4 I__11148 (
            .O(N__47811),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__11147 (
            .O(N__47808),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__11146 (
            .O(N__47805),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__11145 (
            .O(N__47798),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CEMux I__11144 (
            .O(N__47795),
            .I(N__47771));
    CEMux I__11143 (
            .O(N__47794),
            .I(N__47771));
    CEMux I__11142 (
            .O(N__47793),
            .I(N__47771));
    CEMux I__11141 (
            .O(N__47792),
            .I(N__47771));
    CEMux I__11140 (
            .O(N__47791),
            .I(N__47771));
    CEMux I__11139 (
            .O(N__47790),
            .I(N__47771));
    CEMux I__11138 (
            .O(N__47789),
            .I(N__47771));
    CEMux I__11137 (
            .O(N__47788),
            .I(N__47771));
    GlobalMux I__11136 (
            .O(N__47771),
            .I(N__47768));
    gio2CtrlBuf I__11135 (
            .O(N__47768),
            .I(\current_shift_inst.timer_s1.N_161_i_g ));
    InMux I__11134 (
            .O(N__47765),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__11133 (
            .O(N__47762),
            .I(N__47759));
    LocalMux I__11132 (
            .O(N__47759),
            .I(N__47754));
    InMux I__11131 (
            .O(N__47758),
            .I(N__47751));
    InMux I__11130 (
            .O(N__47757),
            .I(N__47748));
    Span4Mux_v I__11129 (
            .O(N__47754),
            .I(N__47745));
    LocalMux I__11128 (
            .O(N__47751),
            .I(N__47742));
    LocalMux I__11127 (
            .O(N__47748),
            .I(N__47739));
    Span4Mux_v I__11126 (
            .O(N__47745),
            .I(N__47736));
    Span12Mux_h I__11125 (
            .O(N__47742),
            .I(N__47731));
    Span12Mux_v I__11124 (
            .O(N__47739),
            .I(N__47731));
    Odrv4 I__11123 (
            .O(N__47736),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv12 I__11122 (
            .O(N__47731),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__11121 (
            .O(N__47726),
            .I(N__47723));
    LocalMux I__11120 (
            .O(N__47723),
            .I(N__47719));
    CascadeMux I__11119 (
            .O(N__47722),
            .I(N__47716));
    Span4Mux_h I__11118 (
            .O(N__47719),
            .I(N__47713));
    InMux I__11117 (
            .O(N__47716),
            .I(N__47709));
    Span4Mux_v I__11116 (
            .O(N__47713),
            .I(N__47706));
    InMux I__11115 (
            .O(N__47712),
            .I(N__47703));
    LocalMux I__11114 (
            .O(N__47709),
            .I(N__47700));
    Odrv4 I__11113 (
            .O(N__47706),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__11112 (
            .O(N__47703),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv12 I__11111 (
            .O(N__47700),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__11110 (
            .O(N__47693),
            .I(bfn_18_23_0_));
    CascadeMux I__11109 (
            .O(N__47690),
            .I(N__47686));
    InMux I__11108 (
            .O(N__47689),
            .I(N__47682));
    InMux I__11107 (
            .O(N__47686),
            .I(N__47679));
    InMux I__11106 (
            .O(N__47685),
            .I(N__47676));
    LocalMux I__11105 (
            .O(N__47682),
            .I(N__47672));
    LocalMux I__11104 (
            .O(N__47679),
            .I(N__47667));
    LocalMux I__11103 (
            .O(N__47676),
            .I(N__47667));
    InMux I__11102 (
            .O(N__47675),
            .I(N__47664));
    Span12Mux_h I__11101 (
            .O(N__47672),
            .I(N__47661));
    Span4Mux_v I__11100 (
            .O(N__47667),
            .I(N__47656));
    LocalMux I__11099 (
            .O(N__47664),
            .I(N__47656));
    Odrv12 I__11098 (
            .O(N__47661),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__11097 (
            .O(N__47656),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__11096 (
            .O(N__47651),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__11095 (
            .O(N__47648),
            .I(N__47645));
    InMux I__11094 (
            .O(N__47645),
            .I(N__47640));
    InMux I__11093 (
            .O(N__47644),
            .I(N__47637));
    InMux I__11092 (
            .O(N__47643),
            .I(N__47634));
    LocalMux I__11091 (
            .O(N__47640),
            .I(N__47631));
    LocalMux I__11090 (
            .O(N__47637),
            .I(N__47628));
    LocalMux I__11089 (
            .O(N__47634),
            .I(N__47625));
    Sp12to4 I__11088 (
            .O(N__47631),
            .I(N__47621));
    Span4Mux_v I__11087 (
            .O(N__47628),
            .I(N__47618));
    Span4Mux_v I__11086 (
            .O(N__47625),
            .I(N__47615));
    InMux I__11085 (
            .O(N__47624),
            .I(N__47612));
    Odrv12 I__11084 (
            .O(N__47621),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__11083 (
            .O(N__47618),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__11082 (
            .O(N__47615),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__11081 (
            .O(N__47612),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__11080 (
            .O(N__47603),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__11079 (
            .O(N__47600),
            .I(N__47596));
    InMux I__11078 (
            .O(N__47599),
            .I(N__47592));
    InMux I__11077 (
            .O(N__47596),
            .I(N__47589));
    InMux I__11076 (
            .O(N__47595),
            .I(N__47586));
    LocalMux I__11075 (
            .O(N__47592),
            .I(N__47581));
    LocalMux I__11074 (
            .O(N__47589),
            .I(N__47581));
    LocalMux I__11073 (
            .O(N__47586),
            .I(N__47578));
    Span4Mux_h I__11072 (
            .O(N__47581),
            .I(N__47574));
    Span4Mux_h I__11071 (
            .O(N__47578),
            .I(N__47571));
    InMux I__11070 (
            .O(N__47577),
            .I(N__47568));
    Odrv4 I__11069 (
            .O(N__47574),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__11068 (
            .O(N__47571),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__11067 (
            .O(N__47568),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__11066 (
            .O(N__47561),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__11065 (
            .O(N__47558),
            .I(N__47555));
    InMux I__11064 (
            .O(N__47555),
            .I(N__47551));
    InMux I__11063 (
            .O(N__47554),
            .I(N__47548));
    LocalMux I__11062 (
            .O(N__47551),
            .I(N__47545));
    LocalMux I__11061 (
            .O(N__47548),
            .I(N__47542));
    Span4Mux_v I__11060 (
            .O(N__47545),
            .I(N__47537));
    Span12Mux_v I__11059 (
            .O(N__47542),
            .I(N__47534));
    InMux I__11058 (
            .O(N__47541),
            .I(N__47531));
    InMux I__11057 (
            .O(N__47540),
            .I(N__47528));
    Odrv4 I__11056 (
            .O(N__47537),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv12 I__11055 (
            .O(N__47534),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__11054 (
            .O(N__47531),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__11053 (
            .O(N__47528),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__11052 (
            .O(N__47519),
            .I(bfn_18_21_0_));
    CascadeMux I__11051 (
            .O(N__47516),
            .I(N__47513));
    InMux I__11050 (
            .O(N__47513),
            .I(N__47509));
    CascadeMux I__11049 (
            .O(N__47512),
            .I(N__47506));
    LocalMux I__11048 (
            .O(N__47509),
            .I(N__47503));
    InMux I__11047 (
            .O(N__47506),
            .I(N__47500));
    Span4Mux_h I__11046 (
            .O(N__47503),
            .I(N__47495));
    LocalMux I__11045 (
            .O(N__47500),
            .I(N__47495));
    Span4Mux_v I__11044 (
            .O(N__47495),
            .I(N__47490));
    InMux I__11043 (
            .O(N__47494),
            .I(N__47487));
    InMux I__11042 (
            .O(N__47493),
            .I(N__47484));
    Odrv4 I__11041 (
            .O(N__47490),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__11040 (
            .O(N__47487),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__11039 (
            .O(N__47484),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__11038 (
            .O(N__47477),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__11037 (
            .O(N__47474),
            .I(N__47470));
    CascadeMux I__11036 (
            .O(N__47473),
            .I(N__47467));
    InMux I__11035 (
            .O(N__47470),
            .I(N__47464));
    InMux I__11034 (
            .O(N__47467),
            .I(N__47461));
    LocalMux I__11033 (
            .O(N__47464),
            .I(N__47455));
    LocalMux I__11032 (
            .O(N__47461),
            .I(N__47455));
    InMux I__11031 (
            .O(N__47460),
            .I(N__47452));
    Span4Mux_v I__11030 (
            .O(N__47455),
            .I(N__47447));
    LocalMux I__11029 (
            .O(N__47452),
            .I(N__47447));
    Span4Mux_h I__11028 (
            .O(N__47447),
            .I(N__47443));
    InMux I__11027 (
            .O(N__47446),
            .I(N__47440));
    Odrv4 I__11026 (
            .O(N__47443),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__11025 (
            .O(N__47440),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__11024 (
            .O(N__47435),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__11023 (
            .O(N__47432),
            .I(N__47428));
    InMux I__11022 (
            .O(N__47431),
            .I(N__47425));
    InMux I__11021 (
            .O(N__47428),
            .I(N__47422));
    LocalMux I__11020 (
            .O(N__47425),
            .I(N__47418));
    LocalMux I__11019 (
            .O(N__47422),
            .I(N__47415));
    InMux I__11018 (
            .O(N__47421),
            .I(N__47412));
    Span4Mux_h I__11017 (
            .O(N__47418),
            .I(N__47409));
    Span4Mux_h I__11016 (
            .O(N__47415),
            .I(N__47405));
    LocalMux I__11015 (
            .O(N__47412),
            .I(N__47402));
    Span4Mux_v I__11014 (
            .O(N__47409),
            .I(N__47399));
    InMux I__11013 (
            .O(N__47408),
            .I(N__47396));
    Odrv4 I__11012 (
            .O(N__47405),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv12 I__11011 (
            .O(N__47402),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__11010 (
            .O(N__47399),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__11009 (
            .O(N__47396),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__11008 (
            .O(N__47387),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__11007 (
            .O(N__47384),
            .I(N__47380));
    InMux I__11006 (
            .O(N__47383),
            .I(N__47377));
    InMux I__11005 (
            .O(N__47380),
            .I(N__47374));
    LocalMux I__11004 (
            .O(N__47377),
            .I(N__47371));
    LocalMux I__11003 (
            .O(N__47374),
            .I(N__47368));
    Span4Mux_h I__11002 (
            .O(N__47371),
            .I(N__47363));
    Span4Mux_v I__11001 (
            .O(N__47368),
            .I(N__47360));
    InMux I__11000 (
            .O(N__47367),
            .I(N__47355));
    InMux I__10999 (
            .O(N__47366),
            .I(N__47355));
    Odrv4 I__10998 (
            .O(N__47363),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__10997 (
            .O(N__47360),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__10996 (
            .O(N__47355),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__10995 (
            .O(N__47348),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__10994 (
            .O(N__47345),
            .I(N__47342));
    InMux I__10993 (
            .O(N__47342),
            .I(N__47337));
    InMux I__10992 (
            .O(N__47341),
            .I(N__47334));
    InMux I__10991 (
            .O(N__47340),
            .I(N__47331));
    LocalMux I__10990 (
            .O(N__47337),
            .I(N__47328));
    LocalMux I__10989 (
            .O(N__47334),
            .I(N__47323));
    LocalMux I__10988 (
            .O(N__47331),
            .I(N__47323));
    Span4Mux_v I__10987 (
            .O(N__47328),
            .I(N__47319));
    Span4Mux_v I__10986 (
            .O(N__47323),
            .I(N__47316));
    InMux I__10985 (
            .O(N__47322),
            .I(N__47313));
    Odrv4 I__10984 (
            .O(N__47319),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__10983 (
            .O(N__47316),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__10982 (
            .O(N__47313),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__10981 (
            .O(N__47306),
            .I(N__47302));
    CascadeMux I__10980 (
            .O(N__47305),
            .I(N__47298));
    LocalMux I__10979 (
            .O(N__47302),
            .I(N__47295));
    InMux I__10978 (
            .O(N__47301),
            .I(N__47292));
    InMux I__10977 (
            .O(N__47298),
            .I(N__47289));
    Span4Mux_v I__10976 (
            .O(N__47295),
            .I(N__47284));
    LocalMux I__10975 (
            .O(N__47292),
            .I(N__47284));
    LocalMux I__10974 (
            .O(N__47289),
            .I(N__47278));
    Span4Mux_v I__10973 (
            .O(N__47284),
            .I(N__47278));
    InMux I__10972 (
            .O(N__47283),
            .I(N__47275));
    Span4Mux_h I__10971 (
            .O(N__47278),
            .I(N__47272));
    LocalMux I__10970 (
            .O(N__47275),
            .I(N__47269));
    Odrv4 I__10969 (
            .O(N__47272),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__10968 (
            .O(N__47269),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__10967 (
            .O(N__47264),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__10966 (
            .O(N__47261),
            .I(N__47257));
    InMux I__10965 (
            .O(N__47260),
            .I(N__47252));
    InMux I__10964 (
            .O(N__47257),
            .I(N__47249));
    InMux I__10963 (
            .O(N__47256),
            .I(N__47244));
    InMux I__10962 (
            .O(N__47255),
            .I(N__47244));
    LocalMux I__10961 (
            .O(N__47252),
            .I(N__47241));
    LocalMux I__10960 (
            .O(N__47249),
            .I(N__47238));
    LocalMux I__10959 (
            .O(N__47244),
            .I(N__47235));
    Span4Mux_h I__10958 (
            .O(N__47241),
            .I(N__47232));
    Span4Mux_v I__10957 (
            .O(N__47238),
            .I(N__47227));
    Span4Mux_h I__10956 (
            .O(N__47235),
            .I(N__47227));
    Odrv4 I__10955 (
            .O(N__47232),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__10954 (
            .O(N__47227),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__10953 (
            .O(N__47222),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__10952 (
            .O(N__47219),
            .I(N__47212));
    InMux I__10951 (
            .O(N__47218),
            .I(N__47212));
    InMux I__10950 (
            .O(N__47217),
            .I(N__47209));
    LocalMux I__10949 (
            .O(N__47212),
            .I(N__47204));
    LocalMux I__10948 (
            .O(N__47209),
            .I(N__47204));
    Span4Mux_h I__10947 (
            .O(N__47204),
            .I(N__47201));
    Span4Mux_v I__10946 (
            .O(N__47201),
            .I(N__47197));
    InMux I__10945 (
            .O(N__47200),
            .I(N__47194));
    Odrv4 I__10944 (
            .O(N__47197),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__10943 (
            .O(N__47194),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__10942 (
            .O(N__47189),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__10941 (
            .O(N__47186),
            .I(N__47183));
    InMux I__10940 (
            .O(N__47183),
            .I(N__47180));
    LocalMux I__10939 (
            .O(N__47180),
            .I(N__47175));
    InMux I__10938 (
            .O(N__47179),
            .I(N__47172));
    InMux I__10937 (
            .O(N__47178),
            .I(N__47169));
    Span4Mux_h I__10936 (
            .O(N__47175),
            .I(N__47164));
    LocalMux I__10935 (
            .O(N__47172),
            .I(N__47164));
    LocalMux I__10934 (
            .O(N__47169),
            .I(N__47160));
    Span4Mux_v I__10933 (
            .O(N__47164),
            .I(N__47157));
    InMux I__10932 (
            .O(N__47163),
            .I(N__47154));
    Odrv12 I__10931 (
            .O(N__47160),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__10930 (
            .O(N__47157),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__10929 (
            .O(N__47154),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__10928 (
            .O(N__47147),
            .I(bfn_18_20_0_));
    CascadeMux I__10927 (
            .O(N__47144),
            .I(N__47141));
    InMux I__10926 (
            .O(N__47141),
            .I(N__47137));
    InMux I__10925 (
            .O(N__47140),
            .I(N__47134));
    LocalMux I__10924 (
            .O(N__47137),
            .I(N__47131));
    LocalMux I__10923 (
            .O(N__47134),
            .I(N__47126));
    Span4Mux_h I__10922 (
            .O(N__47131),
            .I(N__47123));
    InMux I__10921 (
            .O(N__47130),
            .I(N__47118));
    InMux I__10920 (
            .O(N__47129),
            .I(N__47118));
    Span4Mux_h I__10919 (
            .O(N__47126),
            .I(N__47113));
    Span4Mux_v I__10918 (
            .O(N__47123),
            .I(N__47113));
    LocalMux I__10917 (
            .O(N__47118),
            .I(N__47110));
    Odrv4 I__10916 (
            .O(N__47113),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv12 I__10915 (
            .O(N__47110),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10914 (
            .O(N__47105),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__10913 (
            .O(N__47102),
            .I(N__47099));
    InMux I__10912 (
            .O(N__47099),
            .I(N__47095));
    InMux I__10911 (
            .O(N__47098),
            .I(N__47092));
    LocalMux I__10910 (
            .O(N__47095),
            .I(N__47085));
    LocalMux I__10909 (
            .O(N__47092),
            .I(N__47085));
    InMux I__10908 (
            .O(N__47091),
            .I(N__47082));
    InMux I__10907 (
            .O(N__47090),
            .I(N__47079));
    Span4Mux_v I__10906 (
            .O(N__47085),
            .I(N__47076));
    LocalMux I__10905 (
            .O(N__47082),
            .I(N__47073));
    LocalMux I__10904 (
            .O(N__47079),
            .I(N__47070));
    Odrv4 I__10903 (
            .O(N__47076),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv12 I__10902 (
            .O(N__47073),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__10901 (
            .O(N__47070),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__10900 (
            .O(N__47063),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__10899 (
            .O(N__47060),
            .I(N__47057));
    InMux I__10898 (
            .O(N__47057),
            .I(N__47053));
    CascadeMux I__10897 (
            .O(N__47056),
            .I(N__47050));
    LocalMux I__10896 (
            .O(N__47053),
            .I(N__47045));
    InMux I__10895 (
            .O(N__47050),
            .I(N__47042));
    InMux I__10894 (
            .O(N__47049),
            .I(N__47039));
    InMux I__10893 (
            .O(N__47048),
            .I(N__47036));
    Span4Mux_h I__10892 (
            .O(N__47045),
            .I(N__47033));
    LocalMux I__10891 (
            .O(N__47042),
            .I(N__47028));
    LocalMux I__10890 (
            .O(N__47039),
            .I(N__47028));
    LocalMux I__10889 (
            .O(N__47036),
            .I(N__47025));
    Span4Mux_v I__10888 (
            .O(N__47033),
            .I(N__47020));
    Span4Mux_h I__10887 (
            .O(N__47028),
            .I(N__47020));
    Odrv12 I__10886 (
            .O(N__47025),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__10885 (
            .O(N__47020),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__10884 (
            .O(N__47015),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__10883 (
            .O(N__47012),
            .I(N__47008));
    InMux I__10882 (
            .O(N__47011),
            .I(N__47004));
    LocalMux I__10881 (
            .O(N__47008),
            .I(N__47000));
    InMux I__10880 (
            .O(N__47007),
            .I(N__46997));
    LocalMux I__10879 (
            .O(N__47004),
            .I(N__46994));
    InMux I__10878 (
            .O(N__47003),
            .I(N__46991));
    Span4Mux_v I__10877 (
            .O(N__47000),
            .I(N__46988));
    LocalMux I__10876 (
            .O(N__46997),
            .I(N__46985));
    Span4Mux_v I__10875 (
            .O(N__46994),
            .I(N__46980));
    LocalMux I__10874 (
            .O(N__46991),
            .I(N__46980));
    Odrv4 I__10873 (
            .O(N__46988),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv12 I__10872 (
            .O(N__46985),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__10871 (
            .O(N__46980),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__10870 (
            .O(N__46973),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__10869 (
            .O(N__46970),
            .I(N__46967));
    LocalMux I__10868 (
            .O(N__46967),
            .I(N__46964));
    Span4Mux_v I__10867 (
            .O(N__46964),
            .I(N__46961));
    Odrv4 I__10866 (
            .O(N__46961),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__10865 (
            .O(N__46958),
            .I(N__46955));
    LocalMux I__10864 (
            .O(N__46955),
            .I(N__46952));
    Odrv4 I__10863 (
            .O(N__46952),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__10862 (
            .O(N__46949),
            .I(N__46946));
    LocalMux I__10861 (
            .O(N__46946),
            .I(N__46943));
    Odrv4 I__10860 (
            .O(N__46943),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__10859 (
            .O(N__46940),
            .I(N__46937));
    LocalMux I__10858 (
            .O(N__46937),
            .I(N__46934));
    Odrv4 I__10857 (
            .O(N__46934),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    CascadeMux I__10856 (
            .O(N__46931),
            .I(N__46927));
    CascadeMux I__10855 (
            .O(N__46930),
            .I(N__46924));
    InMux I__10854 (
            .O(N__46927),
            .I(N__46921));
    InMux I__10853 (
            .O(N__46924),
            .I(N__46918));
    LocalMux I__10852 (
            .O(N__46921),
            .I(N__46914));
    LocalMux I__10851 (
            .O(N__46918),
            .I(N__46911));
    InMux I__10850 (
            .O(N__46917),
            .I(N__46908));
    Span4Mux_v I__10849 (
            .O(N__46914),
            .I(N__46905));
    Span4Mux_v I__10848 (
            .O(N__46911),
            .I(N__46899));
    LocalMux I__10847 (
            .O(N__46908),
            .I(N__46899));
    Span4Mux_v I__10846 (
            .O(N__46905),
            .I(N__46896));
    InMux I__10845 (
            .O(N__46904),
            .I(N__46893));
    Span4Mux_h I__10844 (
            .O(N__46899),
            .I(N__46890));
    Span4Mux_h I__10843 (
            .O(N__46896),
            .I(N__46885));
    LocalMux I__10842 (
            .O(N__46893),
            .I(N__46885));
    Odrv4 I__10841 (
            .O(N__46890),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__10840 (
            .O(N__46885),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    CascadeMux I__10839 (
            .O(N__46880),
            .I(N__46876));
    CascadeMux I__10838 (
            .O(N__46879),
            .I(N__46873));
    InMux I__10837 (
            .O(N__46876),
            .I(N__46868));
    InMux I__10836 (
            .O(N__46873),
            .I(N__46868));
    LocalMux I__10835 (
            .O(N__46868),
            .I(N__46864));
    InMux I__10834 (
            .O(N__46867),
            .I(N__46861));
    Span4Mux_v I__10833 (
            .O(N__46864),
            .I(N__46856));
    LocalMux I__10832 (
            .O(N__46861),
            .I(N__46856));
    Span4Mux_h I__10831 (
            .O(N__46856),
            .I(N__46852));
    InMux I__10830 (
            .O(N__46855),
            .I(N__46849));
    Odrv4 I__10829 (
            .O(N__46852),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__10828 (
            .O(N__46849),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__10827 (
            .O(N__46844),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__10826 (
            .O(N__46841),
            .I(N__46837));
    CascadeMux I__10825 (
            .O(N__46840),
            .I(N__46834));
    InMux I__10824 (
            .O(N__46837),
            .I(N__46831));
    InMux I__10823 (
            .O(N__46834),
            .I(N__46828));
    LocalMux I__10822 (
            .O(N__46831),
            .I(N__46822));
    LocalMux I__10821 (
            .O(N__46828),
            .I(N__46822));
    InMux I__10820 (
            .O(N__46827),
            .I(N__46819));
    Span4Mux_v I__10819 (
            .O(N__46822),
            .I(N__46815));
    LocalMux I__10818 (
            .O(N__46819),
            .I(N__46812));
    InMux I__10817 (
            .O(N__46818),
            .I(N__46809));
    Span4Mux_v I__10816 (
            .O(N__46815),
            .I(N__46806));
    Span4Mux_h I__10815 (
            .O(N__46812),
            .I(N__46801));
    LocalMux I__10814 (
            .O(N__46809),
            .I(N__46801));
    Odrv4 I__10813 (
            .O(N__46806),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__10812 (
            .O(N__46801),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__10811 (
            .O(N__46796),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__10810 (
            .O(N__46793),
            .I(N__46790));
    InMux I__10809 (
            .O(N__46790),
            .I(N__46786));
    CascadeMux I__10808 (
            .O(N__46789),
            .I(N__46783));
    LocalMux I__10807 (
            .O(N__46786),
            .I(N__46778));
    InMux I__10806 (
            .O(N__46783),
            .I(N__46775));
    InMux I__10805 (
            .O(N__46782),
            .I(N__46772));
    InMux I__10804 (
            .O(N__46781),
            .I(N__46769));
    Span4Mux_v I__10803 (
            .O(N__46778),
            .I(N__46766));
    LocalMux I__10802 (
            .O(N__46775),
            .I(N__46763));
    LocalMux I__10801 (
            .O(N__46772),
            .I(N__46760));
    LocalMux I__10800 (
            .O(N__46769),
            .I(N__46757));
    Span4Mux_v I__10799 (
            .O(N__46766),
            .I(N__46754));
    Span4Mux_v I__10798 (
            .O(N__46763),
            .I(N__46749));
    Span4Mux_h I__10797 (
            .O(N__46760),
            .I(N__46749));
    Span4Mux_v I__10796 (
            .O(N__46757),
            .I(N__46746));
    Odrv4 I__10795 (
            .O(N__46754),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__10794 (
            .O(N__46749),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__10793 (
            .O(N__46746),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__10792 (
            .O(N__46739),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__10791 (
            .O(N__46736),
            .I(N__46732));
    InMux I__10790 (
            .O(N__46735),
            .I(N__46728));
    LocalMux I__10789 (
            .O(N__46732),
            .I(N__46725));
    InMux I__10788 (
            .O(N__46731),
            .I(N__46722));
    LocalMux I__10787 (
            .O(N__46728),
            .I(N__46715));
    Span4Mux_v I__10786 (
            .O(N__46725),
            .I(N__46715));
    LocalMux I__10785 (
            .O(N__46722),
            .I(N__46715));
    Span4Mux_v I__10784 (
            .O(N__46715),
            .I(N__46711));
    InMux I__10783 (
            .O(N__46714),
            .I(N__46708));
    Odrv4 I__10782 (
            .O(N__46711),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__10781 (
            .O(N__46708),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__10780 (
            .O(N__46703),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__10779 (
            .O(N__46700),
            .I(N__46696));
    InMux I__10778 (
            .O(N__46699),
            .I(N__46693));
    InMux I__10777 (
            .O(N__46696),
            .I(N__46690));
    LocalMux I__10776 (
            .O(N__46693),
            .I(N__46687));
    LocalMux I__10775 (
            .O(N__46690),
            .I(N__46681));
    Span4Mux_h I__10774 (
            .O(N__46687),
            .I(N__46681));
    InMux I__10773 (
            .O(N__46686),
            .I(N__46678));
    Odrv4 I__10772 (
            .O(N__46681),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__10771 (
            .O(N__46678),
            .I(\current_shift_inst.un4_control_input1_9 ));
    CascadeMux I__10770 (
            .O(N__46673),
            .I(N__46670));
    InMux I__10769 (
            .O(N__46670),
            .I(N__46667));
    LocalMux I__10768 (
            .O(N__46667),
            .I(N__46664));
    Odrv12 I__10767 (
            .O(N__46664),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    CascadeMux I__10766 (
            .O(N__46661),
            .I(N__46654));
    CascadeMux I__10765 (
            .O(N__46660),
            .I(N__46639));
    CascadeMux I__10764 (
            .O(N__46659),
            .I(N__46633));
    InMux I__10763 (
            .O(N__46658),
            .I(N__46614));
    InMux I__10762 (
            .O(N__46657),
            .I(N__46614));
    InMux I__10761 (
            .O(N__46654),
            .I(N__46614));
    CascadeMux I__10760 (
            .O(N__46653),
            .I(N__46611));
    CascadeMux I__10759 (
            .O(N__46652),
            .I(N__46607));
    CascadeMux I__10758 (
            .O(N__46651),
            .I(N__46584));
    InMux I__10757 (
            .O(N__46650),
            .I(N__46567));
    InMux I__10756 (
            .O(N__46649),
            .I(N__46567));
    InMux I__10755 (
            .O(N__46648),
            .I(N__46567));
    InMux I__10754 (
            .O(N__46647),
            .I(N__46567));
    InMux I__10753 (
            .O(N__46646),
            .I(N__46567));
    InMux I__10752 (
            .O(N__46645),
            .I(N__46567));
    InMux I__10751 (
            .O(N__46644),
            .I(N__46567));
    InMux I__10750 (
            .O(N__46643),
            .I(N__46567));
    InMux I__10749 (
            .O(N__46642),
            .I(N__46543));
    InMux I__10748 (
            .O(N__46639),
            .I(N__46543));
    InMux I__10747 (
            .O(N__46638),
            .I(N__46543));
    InMux I__10746 (
            .O(N__46637),
            .I(N__46543));
    InMux I__10745 (
            .O(N__46636),
            .I(N__46543));
    InMux I__10744 (
            .O(N__46633),
            .I(N__46543));
    InMux I__10743 (
            .O(N__46632),
            .I(N__46543));
    InMux I__10742 (
            .O(N__46631),
            .I(N__46543));
    InMux I__10741 (
            .O(N__46630),
            .I(N__46528));
    InMux I__10740 (
            .O(N__46629),
            .I(N__46528));
    InMux I__10739 (
            .O(N__46628),
            .I(N__46528));
    InMux I__10738 (
            .O(N__46627),
            .I(N__46528));
    InMux I__10737 (
            .O(N__46626),
            .I(N__46528));
    InMux I__10736 (
            .O(N__46625),
            .I(N__46528));
    InMux I__10735 (
            .O(N__46624),
            .I(N__46528));
    CascadeMux I__10734 (
            .O(N__46623),
            .I(N__46520));
    CascadeMux I__10733 (
            .O(N__46622),
            .I(N__46517));
    CascadeMux I__10732 (
            .O(N__46621),
            .I(N__46514));
    LocalMux I__10731 (
            .O(N__46614),
            .I(N__46501));
    InMux I__10730 (
            .O(N__46611),
            .I(N__46484));
    InMux I__10729 (
            .O(N__46610),
            .I(N__46484));
    InMux I__10728 (
            .O(N__46607),
            .I(N__46484));
    InMux I__10727 (
            .O(N__46606),
            .I(N__46484));
    InMux I__10726 (
            .O(N__46605),
            .I(N__46484));
    InMux I__10725 (
            .O(N__46604),
            .I(N__46484));
    InMux I__10724 (
            .O(N__46603),
            .I(N__46484));
    InMux I__10723 (
            .O(N__46602),
            .I(N__46484));
    InMux I__10722 (
            .O(N__46601),
            .I(N__46481));
    CascadeMux I__10721 (
            .O(N__46600),
            .I(N__46478));
    CascadeMux I__10720 (
            .O(N__46599),
            .I(N__46474));
    CascadeMux I__10719 (
            .O(N__46598),
            .I(N__46470));
    CascadeMux I__10718 (
            .O(N__46597),
            .I(N__46466));
    CascadeMux I__10717 (
            .O(N__46596),
            .I(N__46463));
    CascadeMux I__10716 (
            .O(N__46595),
            .I(N__46459));
    CascadeMux I__10715 (
            .O(N__46594),
            .I(N__46455));
    CascadeMux I__10714 (
            .O(N__46593),
            .I(N__46451));
    CascadeMux I__10713 (
            .O(N__46592),
            .I(N__46435));
    CascadeMux I__10712 (
            .O(N__46591),
            .I(N__46431));
    CascadeMux I__10711 (
            .O(N__46590),
            .I(N__46427));
    InMux I__10710 (
            .O(N__46589),
            .I(N__46420));
    InMux I__10709 (
            .O(N__46588),
            .I(N__46420));
    InMux I__10708 (
            .O(N__46587),
            .I(N__46420));
    InMux I__10707 (
            .O(N__46584),
            .I(N__46417));
    LocalMux I__10706 (
            .O(N__46567),
            .I(N__46414));
    InMux I__10705 (
            .O(N__46566),
            .I(N__46399));
    InMux I__10704 (
            .O(N__46565),
            .I(N__46399));
    InMux I__10703 (
            .O(N__46564),
            .I(N__46399));
    InMux I__10702 (
            .O(N__46563),
            .I(N__46399));
    InMux I__10701 (
            .O(N__46562),
            .I(N__46399));
    InMux I__10700 (
            .O(N__46561),
            .I(N__46399));
    InMux I__10699 (
            .O(N__46560),
            .I(N__46399));
    LocalMux I__10698 (
            .O(N__46543),
            .I(N__46394));
    LocalMux I__10697 (
            .O(N__46528),
            .I(N__46394));
    InMux I__10696 (
            .O(N__46527),
            .I(N__46389));
    InMux I__10695 (
            .O(N__46526),
            .I(N__46389));
    InMux I__10694 (
            .O(N__46525),
            .I(N__46378));
    InMux I__10693 (
            .O(N__46524),
            .I(N__46378));
    InMux I__10692 (
            .O(N__46523),
            .I(N__46378));
    InMux I__10691 (
            .O(N__46520),
            .I(N__46378));
    InMux I__10690 (
            .O(N__46517),
            .I(N__46378));
    InMux I__10689 (
            .O(N__46514),
            .I(N__46368));
    InMux I__10688 (
            .O(N__46513),
            .I(N__46368));
    InMux I__10687 (
            .O(N__46512),
            .I(N__46368));
    CascadeMux I__10686 (
            .O(N__46511),
            .I(N__46364));
    CascadeMux I__10685 (
            .O(N__46510),
            .I(N__46360));
    CascadeMux I__10684 (
            .O(N__46509),
            .I(N__46356));
    CascadeMux I__10683 (
            .O(N__46508),
            .I(N__46352));
    CascadeMux I__10682 (
            .O(N__46507),
            .I(N__46349));
    CascadeMux I__10681 (
            .O(N__46506),
            .I(N__46345));
    CascadeMux I__10680 (
            .O(N__46505),
            .I(N__46341));
    CascadeMux I__10679 (
            .O(N__46504),
            .I(N__46337));
    Span4Mux_v I__10678 (
            .O(N__46501),
            .I(N__46333));
    LocalMux I__10677 (
            .O(N__46484),
            .I(N__46328));
    LocalMux I__10676 (
            .O(N__46481),
            .I(N__46328));
    InMux I__10675 (
            .O(N__46478),
            .I(N__46313));
    InMux I__10674 (
            .O(N__46477),
            .I(N__46313));
    InMux I__10673 (
            .O(N__46474),
            .I(N__46313));
    InMux I__10672 (
            .O(N__46473),
            .I(N__46313));
    InMux I__10671 (
            .O(N__46470),
            .I(N__46313));
    InMux I__10670 (
            .O(N__46469),
            .I(N__46313));
    InMux I__10669 (
            .O(N__46466),
            .I(N__46313));
    InMux I__10668 (
            .O(N__46463),
            .I(N__46296));
    InMux I__10667 (
            .O(N__46462),
            .I(N__46296));
    InMux I__10666 (
            .O(N__46459),
            .I(N__46296));
    InMux I__10665 (
            .O(N__46458),
            .I(N__46296));
    InMux I__10664 (
            .O(N__46455),
            .I(N__46296));
    InMux I__10663 (
            .O(N__46454),
            .I(N__46296));
    InMux I__10662 (
            .O(N__46451),
            .I(N__46296));
    InMux I__10661 (
            .O(N__46450),
            .I(N__46296));
    CascadeMux I__10660 (
            .O(N__46449),
            .I(N__46293));
    CascadeMux I__10659 (
            .O(N__46448),
            .I(N__46289));
    CascadeMux I__10658 (
            .O(N__46447),
            .I(N__46285));
    CascadeMux I__10657 (
            .O(N__46446),
            .I(N__46281));
    CascadeMux I__10656 (
            .O(N__46445),
            .I(N__46277));
    CascadeMux I__10655 (
            .O(N__46444),
            .I(N__46273));
    CascadeMux I__10654 (
            .O(N__46443),
            .I(N__46269));
    CascadeMux I__10653 (
            .O(N__46442),
            .I(N__46265));
    CascadeMux I__10652 (
            .O(N__46441),
            .I(N__46261));
    CascadeMux I__10651 (
            .O(N__46440),
            .I(N__46257));
    CascadeMux I__10650 (
            .O(N__46439),
            .I(N__46253));
    InMux I__10649 (
            .O(N__46438),
            .I(N__46239));
    InMux I__10648 (
            .O(N__46435),
            .I(N__46239));
    InMux I__10647 (
            .O(N__46434),
            .I(N__46239));
    InMux I__10646 (
            .O(N__46431),
            .I(N__46239));
    InMux I__10645 (
            .O(N__46430),
            .I(N__46239));
    InMux I__10644 (
            .O(N__46427),
            .I(N__46239));
    LocalMux I__10643 (
            .O(N__46420),
            .I(N__46236));
    LocalMux I__10642 (
            .O(N__46417),
            .I(N__46229));
    Span12Mux_s11_h I__10641 (
            .O(N__46414),
            .I(N__46229));
    LocalMux I__10640 (
            .O(N__46399),
            .I(N__46229));
    Span4Mux_v I__10639 (
            .O(N__46394),
            .I(N__46222));
    LocalMux I__10638 (
            .O(N__46389),
            .I(N__46222));
    LocalMux I__10637 (
            .O(N__46378),
            .I(N__46222));
    InMux I__10636 (
            .O(N__46377),
            .I(N__46215));
    InMux I__10635 (
            .O(N__46376),
            .I(N__46215));
    InMux I__10634 (
            .O(N__46375),
            .I(N__46215));
    LocalMux I__10633 (
            .O(N__46368),
            .I(N__46212));
    InMux I__10632 (
            .O(N__46367),
            .I(N__46195));
    InMux I__10631 (
            .O(N__46364),
            .I(N__46195));
    InMux I__10630 (
            .O(N__46363),
            .I(N__46195));
    InMux I__10629 (
            .O(N__46360),
            .I(N__46195));
    InMux I__10628 (
            .O(N__46359),
            .I(N__46195));
    InMux I__10627 (
            .O(N__46356),
            .I(N__46195));
    InMux I__10626 (
            .O(N__46355),
            .I(N__46195));
    InMux I__10625 (
            .O(N__46352),
            .I(N__46195));
    InMux I__10624 (
            .O(N__46349),
            .I(N__46178));
    InMux I__10623 (
            .O(N__46348),
            .I(N__46178));
    InMux I__10622 (
            .O(N__46345),
            .I(N__46178));
    InMux I__10621 (
            .O(N__46344),
            .I(N__46178));
    InMux I__10620 (
            .O(N__46341),
            .I(N__46178));
    InMux I__10619 (
            .O(N__46340),
            .I(N__46178));
    InMux I__10618 (
            .O(N__46337),
            .I(N__46178));
    InMux I__10617 (
            .O(N__46336),
            .I(N__46178));
    Span4Mux_h I__10616 (
            .O(N__46333),
            .I(N__46169));
    Span4Mux_h I__10615 (
            .O(N__46328),
            .I(N__46169));
    LocalMux I__10614 (
            .O(N__46313),
            .I(N__46169));
    LocalMux I__10613 (
            .O(N__46296),
            .I(N__46169));
    InMux I__10612 (
            .O(N__46293),
            .I(N__46152));
    InMux I__10611 (
            .O(N__46292),
            .I(N__46152));
    InMux I__10610 (
            .O(N__46289),
            .I(N__46152));
    InMux I__10609 (
            .O(N__46288),
            .I(N__46152));
    InMux I__10608 (
            .O(N__46285),
            .I(N__46152));
    InMux I__10607 (
            .O(N__46284),
            .I(N__46152));
    InMux I__10606 (
            .O(N__46281),
            .I(N__46152));
    InMux I__10605 (
            .O(N__46280),
            .I(N__46152));
    InMux I__10604 (
            .O(N__46277),
            .I(N__46135));
    InMux I__10603 (
            .O(N__46276),
            .I(N__46135));
    InMux I__10602 (
            .O(N__46273),
            .I(N__46135));
    InMux I__10601 (
            .O(N__46272),
            .I(N__46135));
    InMux I__10600 (
            .O(N__46269),
            .I(N__46135));
    InMux I__10599 (
            .O(N__46268),
            .I(N__46135));
    InMux I__10598 (
            .O(N__46265),
            .I(N__46135));
    InMux I__10597 (
            .O(N__46264),
            .I(N__46135));
    InMux I__10596 (
            .O(N__46261),
            .I(N__46122));
    InMux I__10595 (
            .O(N__46260),
            .I(N__46122));
    InMux I__10594 (
            .O(N__46257),
            .I(N__46122));
    InMux I__10593 (
            .O(N__46256),
            .I(N__46122));
    InMux I__10592 (
            .O(N__46253),
            .I(N__46122));
    InMux I__10591 (
            .O(N__46252),
            .I(N__46122));
    LocalMux I__10590 (
            .O(N__46239),
            .I(N__46119));
    Odrv12 I__10589 (
            .O(N__46236),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__10588 (
            .O(N__46229),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10587 (
            .O(N__46222),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10586 (
            .O(N__46215),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10585 (
            .O(N__46212),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10584 (
            .O(N__46195),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10583 (
            .O(N__46178),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10582 (
            .O(N__46169),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10581 (
            .O(N__46152),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10580 (
            .O(N__46135),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10579 (
            .O(N__46122),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10578 (
            .O(N__46119),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__10577 (
            .O(N__46094),
            .I(N__46089));
    InMux I__10576 (
            .O(N__46093),
            .I(N__46086));
    InMux I__10575 (
            .O(N__46092),
            .I(N__46083));
    LocalMux I__10574 (
            .O(N__46089),
            .I(N__46080));
    LocalMux I__10573 (
            .O(N__46086),
            .I(N__46077));
    LocalMux I__10572 (
            .O(N__46083),
            .I(N__46074));
    Span4Mux_h I__10571 (
            .O(N__46080),
            .I(N__46071));
    Span4Mux_h I__10570 (
            .O(N__46077),
            .I(N__46068));
    Span4Mux_h I__10569 (
            .O(N__46074),
            .I(N__46065));
    Odrv4 I__10568 (
            .O(N__46071),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__10567 (
            .O(N__46068),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__10566 (
            .O(N__46065),
            .I(\current_shift_inst.un4_control_input1_11 ));
    CascadeMux I__10565 (
            .O(N__46058),
            .I(N__46055));
    InMux I__10564 (
            .O(N__46055),
            .I(N__46052));
    LocalMux I__10563 (
            .O(N__46052),
            .I(N__46049));
    Odrv12 I__10562 (
            .O(N__46049),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    InMux I__10561 (
            .O(N__46046),
            .I(N__46042));
    InMux I__10560 (
            .O(N__46045),
            .I(N__46038));
    LocalMux I__10559 (
            .O(N__46042),
            .I(N__46035));
    InMux I__10558 (
            .O(N__46041),
            .I(N__46032));
    LocalMux I__10557 (
            .O(N__46038),
            .I(N__46029));
    Span4Mux_h I__10556 (
            .O(N__46035),
            .I(N__46026));
    LocalMux I__10555 (
            .O(N__46032),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv12 I__10554 (
            .O(N__46029),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__10553 (
            .O(N__46026),
            .I(\current_shift_inst.un4_control_input1_14 ));
    CascadeMux I__10552 (
            .O(N__46019),
            .I(N__46016));
    InMux I__10551 (
            .O(N__46016),
            .I(N__46013));
    LocalMux I__10550 (
            .O(N__46013),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__10549 (
            .O(N__46010),
            .I(N__45996));
    CascadeMux I__10548 (
            .O(N__46009),
            .I(N__45988));
    InMux I__10547 (
            .O(N__46008),
            .I(N__45975));
    InMux I__10546 (
            .O(N__46007),
            .I(N__45975));
    InMux I__10545 (
            .O(N__46006),
            .I(N__45975));
    InMux I__10544 (
            .O(N__46005),
            .I(N__45975));
    InMux I__10543 (
            .O(N__46004),
            .I(N__45966));
    InMux I__10542 (
            .O(N__46003),
            .I(N__45966));
    InMux I__10541 (
            .O(N__46002),
            .I(N__45966));
    InMux I__10540 (
            .O(N__46001),
            .I(N__45966));
    InMux I__10539 (
            .O(N__46000),
            .I(N__45963));
    InMux I__10538 (
            .O(N__45999),
            .I(N__45952));
    LocalMux I__10537 (
            .O(N__45996),
            .I(N__45949));
    InMux I__10536 (
            .O(N__45995),
            .I(N__45944));
    InMux I__10535 (
            .O(N__45994),
            .I(N__45944));
    InMux I__10534 (
            .O(N__45993),
            .I(N__45937));
    InMux I__10533 (
            .O(N__45992),
            .I(N__45937));
    InMux I__10532 (
            .O(N__45991),
            .I(N__45937));
    InMux I__10531 (
            .O(N__45988),
            .I(N__45926));
    InMux I__10530 (
            .O(N__45987),
            .I(N__45926));
    InMux I__10529 (
            .O(N__45986),
            .I(N__45926));
    InMux I__10528 (
            .O(N__45985),
            .I(N__45926));
    InMux I__10527 (
            .O(N__45984),
            .I(N__45926));
    LocalMux I__10526 (
            .O(N__45975),
            .I(N__45919));
    LocalMux I__10525 (
            .O(N__45966),
            .I(N__45919));
    LocalMux I__10524 (
            .O(N__45963),
            .I(N__45919));
    InMux I__10523 (
            .O(N__45962),
            .I(N__45900));
    InMux I__10522 (
            .O(N__45961),
            .I(N__45900));
    InMux I__10521 (
            .O(N__45960),
            .I(N__45900));
    InMux I__10520 (
            .O(N__45959),
            .I(N__45891));
    InMux I__10519 (
            .O(N__45958),
            .I(N__45891));
    InMux I__10518 (
            .O(N__45957),
            .I(N__45891));
    InMux I__10517 (
            .O(N__45956),
            .I(N__45891));
    InMux I__10516 (
            .O(N__45955),
            .I(N__45888));
    LocalMux I__10515 (
            .O(N__45952),
            .I(N__45856));
    Span4Mux_h I__10514 (
            .O(N__45949),
            .I(N__45856));
    LocalMux I__10513 (
            .O(N__45944),
            .I(N__45856));
    LocalMux I__10512 (
            .O(N__45937),
            .I(N__45856));
    LocalMux I__10511 (
            .O(N__45926),
            .I(N__45856));
    Span4Mux_v I__10510 (
            .O(N__45919),
            .I(N__45856));
    InMux I__10509 (
            .O(N__45918),
            .I(N__45839));
    InMux I__10508 (
            .O(N__45917),
            .I(N__45839));
    InMux I__10507 (
            .O(N__45916),
            .I(N__45839));
    InMux I__10506 (
            .O(N__45915),
            .I(N__45839));
    InMux I__10505 (
            .O(N__45914),
            .I(N__45839));
    InMux I__10504 (
            .O(N__45913),
            .I(N__45839));
    InMux I__10503 (
            .O(N__45912),
            .I(N__45839));
    InMux I__10502 (
            .O(N__45911),
            .I(N__45839));
    CascadeMux I__10501 (
            .O(N__45910),
            .I(N__45827));
    InMux I__10500 (
            .O(N__45909),
            .I(N__45819));
    InMux I__10499 (
            .O(N__45908),
            .I(N__45819));
    InMux I__10498 (
            .O(N__45907),
            .I(N__45819));
    LocalMux I__10497 (
            .O(N__45900),
            .I(N__45814));
    LocalMux I__10496 (
            .O(N__45891),
            .I(N__45814));
    LocalMux I__10495 (
            .O(N__45888),
            .I(N__45810));
    InMux I__10494 (
            .O(N__45887),
            .I(N__45795));
    InMux I__10493 (
            .O(N__45886),
            .I(N__45795));
    InMux I__10492 (
            .O(N__45885),
            .I(N__45795));
    InMux I__10491 (
            .O(N__45884),
            .I(N__45795));
    InMux I__10490 (
            .O(N__45883),
            .I(N__45795));
    InMux I__10489 (
            .O(N__45882),
            .I(N__45795));
    InMux I__10488 (
            .O(N__45881),
            .I(N__45795));
    InMux I__10487 (
            .O(N__45880),
            .I(N__45780));
    InMux I__10486 (
            .O(N__45879),
            .I(N__45780));
    InMux I__10485 (
            .O(N__45878),
            .I(N__45780));
    InMux I__10484 (
            .O(N__45877),
            .I(N__45780));
    InMux I__10483 (
            .O(N__45876),
            .I(N__45780));
    InMux I__10482 (
            .O(N__45875),
            .I(N__45780));
    InMux I__10481 (
            .O(N__45874),
            .I(N__45780));
    InMux I__10480 (
            .O(N__45873),
            .I(N__45775));
    InMux I__10479 (
            .O(N__45872),
            .I(N__45775));
    InMux I__10478 (
            .O(N__45871),
            .I(N__45768));
    InMux I__10477 (
            .O(N__45870),
            .I(N__45768));
    InMux I__10476 (
            .O(N__45869),
            .I(N__45768));
    Span4Mux_v I__10475 (
            .O(N__45856),
            .I(N__45763));
    LocalMux I__10474 (
            .O(N__45839),
            .I(N__45763));
    InMux I__10473 (
            .O(N__45838),
            .I(N__45752));
    InMux I__10472 (
            .O(N__45837),
            .I(N__45752));
    InMux I__10471 (
            .O(N__45836),
            .I(N__45752));
    InMux I__10470 (
            .O(N__45835),
            .I(N__45752));
    InMux I__10469 (
            .O(N__45834),
            .I(N__45752));
    InMux I__10468 (
            .O(N__45833),
            .I(N__45745));
    InMux I__10467 (
            .O(N__45832),
            .I(N__45745));
    InMux I__10466 (
            .O(N__45831),
            .I(N__45745));
    InMux I__10465 (
            .O(N__45830),
            .I(N__45738));
    InMux I__10464 (
            .O(N__45827),
            .I(N__45738));
    InMux I__10463 (
            .O(N__45826),
            .I(N__45738));
    LocalMux I__10462 (
            .O(N__45819),
            .I(N__45733));
    Span4Mux_v I__10461 (
            .O(N__45814),
            .I(N__45733));
    InMux I__10460 (
            .O(N__45813),
            .I(N__45730));
    Span12Mux_s11_v I__10459 (
            .O(N__45810),
            .I(N__45719));
    LocalMux I__10458 (
            .O(N__45795),
            .I(N__45719));
    LocalMux I__10457 (
            .O(N__45780),
            .I(N__45719));
    LocalMux I__10456 (
            .O(N__45775),
            .I(N__45719));
    LocalMux I__10455 (
            .O(N__45768),
            .I(N__45719));
    Span4Mux_v I__10454 (
            .O(N__45763),
            .I(N__45716));
    LocalMux I__10453 (
            .O(N__45752),
            .I(N__45705));
    LocalMux I__10452 (
            .O(N__45745),
            .I(N__45705));
    LocalMux I__10451 (
            .O(N__45738),
            .I(N__45705));
    Sp12to4 I__10450 (
            .O(N__45733),
            .I(N__45705));
    LocalMux I__10449 (
            .O(N__45730),
            .I(N__45705));
    Span12Mux_s11_h I__10448 (
            .O(N__45719),
            .I(N__45702));
    Odrv4 I__10447 (
            .O(N__45716),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__10446 (
            .O(N__45705),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__10445 (
            .O(N__45702),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__10444 (
            .O(N__45695),
            .I(N__45692));
    LocalMux I__10443 (
            .O(N__45692),
            .I(N__45689));
    Odrv4 I__10442 (
            .O(N__45689),
            .I(\current_shift_inst.un4_control_input1_1 ));
    InMux I__10441 (
            .O(N__45686),
            .I(N__45682));
    InMux I__10440 (
            .O(N__45685),
            .I(N__45679));
    LocalMux I__10439 (
            .O(N__45682),
            .I(N__45676));
    LocalMux I__10438 (
            .O(N__45679),
            .I(N__45673));
    Span4Mux_h I__10437 (
            .O(N__45676),
            .I(N__45668));
    Span4Mux_h I__10436 (
            .O(N__45673),
            .I(N__45665));
    InMux I__10435 (
            .O(N__45672),
            .I(N__45660));
    InMux I__10434 (
            .O(N__45671),
            .I(N__45660));
    Odrv4 I__10433 (
            .O(N__45668),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    Odrv4 I__10432 (
            .O(N__45665),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__10431 (
            .O(N__45660),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__10430 (
            .O(N__45653),
            .I(N__45650));
    InMux I__10429 (
            .O(N__45650),
            .I(N__45647));
    LocalMux I__10428 (
            .O(N__45647),
            .I(N__45644));
    Span4Mux_h I__10427 (
            .O(N__45644),
            .I(N__45641));
    Odrv4 I__10426 (
            .O(N__45641),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__10425 (
            .O(N__45638),
            .I(N__45634));
    InMux I__10424 (
            .O(N__45637),
            .I(N__45631));
    InMux I__10423 (
            .O(N__45634),
            .I(N__45627));
    LocalMux I__10422 (
            .O(N__45631),
            .I(N__45624));
    InMux I__10421 (
            .O(N__45630),
            .I(N__45621));
    LocalMux I__10420 (
            .O(N__45627),
            .I(N__45618));
    Span4Mux_h I__10419 (
            .O(N__45624),
            .I(N__45615));
    LocalMux I__10418 (
            .O(N__45621),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv12 I__10417 (
            .O(N__45618),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__10416 (
            .O(N__45615),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__10415 (
            .O(N__45608),
            .I(N__45605));
    LocalMux I__10414 (
            .O(N__45605),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    InMux I__10413 (
            .O(N__45602),
            .I(N__45599));
    LocalMux I__10412 (
            .O(N__45599),
            .I(N__45596));
    Odrv4 I__10411 (
            .O(N__45596),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__10410 (
            .O(N__45593),
            .I(N__45580));
    InMux I__10409 (
            .O(N__45592),
            .I(N__45580));
    InMux I__10408 (
            .O(N__45591),
            .I(N__45573));
    InMux I__10407 (
            .O(N__45590),
            .I(N__45573));
    InMux I__10406 (
            .O(N__45589),
            .I(N__45573));
    InMux I__10405 (
            .O(N__45588),
            .I(N__45569));
    InMux I__10404 (
            .O(N__45587),
            .I(N__45566));
    InMux I__10403 (
            .O(N__45586),
            .I(N__45561));
    InMux I__10402 (
            .O(N__45585),
            .I(N__45561));
    LocalMux I__10401 (
            .O(N__45580),
            .I(N__45556));
    LocalMux I__10400 (
            .O(N__45573),
            .I(N__45556));
    InMux I__10399 (
            .O(N__45572),
            .I(N__45553));
    LocalMux I__10398 (
            .O(N__45569),
            .I(N__45542));
    LocalMux I__10397 (
            .O(N__45566),
            .I(N__45542));
    LocalMux I__10396 (
            .O(N__45561),
            .I(N__45542));
    Span4Mux_v I__10395 (
            .O(N__45556),
            .I(N__45537));
    LocalMux I__10394 (
            .O(N__45553),
            .I(N__45537));
    InMux I__10393 (
            .O(N__45552),
            .I(N__45528));
    InMux I__10392 (
            .O(N__45551),
            .I(N__45528));
    InMux I__10391 (
            .O(N__45550),
            .I(N__45528));
    InMux I__10390 (
            .O(N__45549),
            .I(N__45528));
    Span4Mux_v I__10389 (
            .O(N__45542),
            .I(N__45514));
    Span4Mux_v I__10388 (
            .O(N__45537),
            .I(N__45509));
    LocalMux I__10387 (
            .O(N__45528),
            .I(N__45509));
    InMux I__10386 (
            .O(N__45527),
            .I(N__45492));
    InMux I__10385 (
            .O(N__45526),
            .I(N__45492));
    InMux I__10384 (
            .O(N__45525),
            .I(N__45492));
    InMux I__10383 (
            .O(N__45524),
            .I(N__45492));
    InMux I__10382 (
            .O(N__45523),
            .I(N__45492));
    InMux I__10381 (
            .O(N__45522),
            .I(N__45492));
    InMux I__10380 (
            .O(N__45521),
            .I(N__45492));
    InMux I__10379 (
            .O(N__45520),
            .I(N__45492));
    InMux I__10378 (
            .O(N__45519),
            .I(N__45489));
    InMux I__10377 (
            .O(N__45518),
            .I(N__45484));
    InMux I__10376 (
            .O(N__45517),
            .I(N__45484));
    Odrv4 I__10375 (
            .O(N__45514),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__10374 (
            .O(N__45509),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10373 (
            .O(N__45492),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10372 (
            .O(N__45489),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10371 (
            .O(N__45484),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__10370 (
            .O(N__45473),
            .I(N__45469));
    InMux I__10369 (
            .O(N__45472),
            .I(N__45466));
    LocalMux I__10368 (
            .O(N__45469),
            .I(N__45462));
    LocalMux I__10367 (
            .O(N__45466),
            .I(N__45459));
    InMux I__10366 (
            .O(N__45465),
            .I(N__45456));
    Span4Mux_h I__10365 (
            .O(N__45462),
            .I(N__45451));
    Span4Mux_v I__10364 (
            .O(N__45459),
            .I(N__45451));
    LocalMux I__10363 (
            .O(N__45456),
            .I(\current_shift_inst.un4_control_input1_21 ));
    Odrv4 I__10362 (
            .O(N__45451),
            .I(\current_shift_inst.un4_control_input1_21 ));
    CascadeMux I__10361 (
            .O(N__45446),
            .I(N__45443));
    InMux I__10360 (
            .O(N__45443),
            .I(N__45440));
    LocalMux I__10359 (
            .O(N__45440),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__10358 (
            .O(N__45437),
            .I(N__45434));
    LocalMux I__10357 (
            .O(N__45434),
            .I(N__45431));
    Odrv4 I__10356 (
            .O(N__45431),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    CascadeMux I__10355 (
            .O(N__45428),
            .I(N__45425));
    InMux I__10354 (
            .O(N__45425),
            .I(N__45422));
    LocalMux I__10353 (
            .O(N__45422),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__10352 (
            .O(N__45419),
            .I(N__45416));
    InMux I__10351 (
            .O(N__45416),
            .I(N__45412));
    CascadeMux I__10350 (
            .O(N__45415),
            .I(N__45409));
    LocalMux I__10349 (
            .O(N__45412),
            .I(N__45405));
    InMux I__10348 (
            .O(N__45409),
            .I(N__45402));
    InMux I__10347 (
            .O(N__45408),
            .I(N__45399));
    Span4Mux_h I__10346 (
            .O(N__45405),
            .I(N__45394));
    LocalMux I__10345 (
            .O(N__45402),
            .I(N__45394));
    LocalMux I__10344 (
            .O(N__45399),
            .I(N__45391));
    Span4Mux_v I__10343 (
            .O(N__45394),
            .I(N__45388));
    Odrv4 I__10342 (
            .O(N__45391),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__10341 (
            .O(N__45388),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__10340 (
            .O(N__45383),
            .I(N__45380));
    InMux I__10339 (
            .O(N__45380),
            .I(N__45377));
    LocalMux I__10338 (
            .O(N__45377),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__10337 (
            .O(N__45374),
            .I(N__45371));
    LocalMux I__10336 (
            .O(N__45371),
            .I(N__45368));
    Span4Mux_h I__10335 (
            .O(N__45368),
            .I(N__45363));
    InMux I__10334 (
            .O(N__45367),
            .I(N__45360));
    InMux I__10333 (
            .O(N__45366),
            .I(N__45357));
    Odrv4 I__10332 (
            .O(N__45363),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__10331 (
            .O(N__45360),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__10330 (
            .O(N__45357),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__10329 (
            .O(N__45350),
            .I(N__45347));
    LocalMux I__10328 (
            .O(N__45347),
            .I(N__45344));
    Odrv4 I__10327 (
            .O(N__45344),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    CascadeMux I__10326 (
            .O(N__45341),
            .I(N__45338));
    InMux I__10325 (
            .O(N__45338),
            .I(N__45335));
    LocalMux I__10324 (
            .O(N__45335),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__10323 (
            .O(N__45332),
            .I(N__45328));
    InMux I__10322 (
            .O(N__45331),
            .I(N__45322));
    InMux I__10321 (
            .O(N__45328),
            .I(N__45322));
    InMux I__10320 (
            .O(N__45327),
            .I(N__45319));
    LocalMux I__10319 (
            .O(N__45322),
            .I(N__45316));
    LocalMux I__10318 (
            .O(N__45319),
            .I(N__45313));
    Span4Mux_h I__10317 (
            .O(N__45316),
            .I(N__45310));
    Span4Mux_h I__10316 (
            .O(N__45313),
            .I(N__45307));
    Odrv4 I__10315 (
            .O(N__45310),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__10314 (
            .O(N__45307),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__10313 (
            .O(N__45302),
            .I(N__45299));
    InMux I__10312 (
            .O(N__45299),
            .I(N__45296));
    LocalMux I__10311 (
            .O(N__45296),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    CascadeMux I__10310 (
            .O(N__45293),
            .I(N__45290));
    InMux I__10309 (
            .O(N__45290),
            .I(N__45287));
    LocalMux I__10308 (
            .O(N__45287),
            .I(N__45282));
    InMux I__10307 (
            .O(N__45286),
            .I(N__45279));
    InMux I__10306 (
            .O(N__45285),
            .I(N__45276));
    Span4Mux_h I__10305 (
            .O(N__45282),
            .I(N__45271));
    LocalMux I__10304 (
            .O(N__45279),
            .I(N__45271));
    LocalMux I__10303 (
            .O(N__45276),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__10302 (
            .O(N__45271),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__10301 (
            .O(N__45266),
            .I(N__45263));
    LocalMux I__10300 (
            .O(N__45263),
            .I(N__45260));
    Odrv4 I__10299 (
            .O(N__45260),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    CascadeMux I__10298 (
            .O(N__45257),
            .I(N__45254));
    InMux I__10297 (
            .O(N__45254),
            .I(N__45251));
    LocalMux I__10296 (
            .O(N__45251),
            .I(N__45246));
    InMux I__10295 (
            .O(N__45250),
            .I(N__45243));
    InMux I__10294 (
            .O(N__45249),
            .I(N__45240));
    Span4Mux_v I__10293 (
            .O(N__45246),
            .I(N__45235));
    LocalMux I__10292 (
            .O(N__45243),
            .I(N__45235));
    LocalMux I__10291 (
            .O(N__45240),
            .I(N__45232));
    Span4Mux_h I__10290 (
            .O(N__45235),
            .I(N__45229));
    Odrv4 I__10289 (
            .O(N__45232),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__10288 (
            .O(N__45229),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__10287 (
            .O(N__45224),
            .I(N__45221));
    InMux I__10286 (
            .O(N__45221),
            .I(N__45218));
    LocalMux I__10285 (
            .O(N__45218),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__10284 (
            .O(N__45215),
            .I(N__45212));
    InMux I__10283 (
            .O(N__45212),
            .I(N__45207));
    InMux I__10282 (
            .O(N__45211),
            .I(N__45204));
    InMux I__10281 (
            .O(N__45210),
            .I(N__45201));
    LocalMux I__10280 (
            .O(N__45207),
            .I(N__45198));
    LocalMux I__10279 (
            .O(N__45204),
            .I(N__45195));
    LocalMux I__10278 (
            .O(N__45201),
            .I(N__45192));
    Span4Mux_v I__10277 (
            .O(N__45198),
            .I(N__45187));
    Span4Mux_h I__10276 (
            .O(N__45195),
            .I(N__45187));
    Span4Mux_h I__10275 (
            .O(N__45192),
            .I(N__45184));
    Odrv4 I__10274 (
            .O(N__45187),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__10273 (
            .O(N__45184),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__10272 (
            .O(N__45179),
            .I(N__45176));
    LocalMux I__10271 (
            .O(N__45176),
            .I(N__45173));
    Odrv12 I__10270 (
            .O(N__45173),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__10269 (
            .O(N__45170),
            .I(N__45165));
    InMux I__10268 (
            .O(N__45169),
            .I(N__45162));
    InMux I__10267 (
            .O(N__45168),
            .I(N__45159));
    LocalMux I__10266 (
            .O(N__45165),
            .I(N__45156));
    LocalMux I__10265 (
            .O(N__45162),
            .I(N__45153));
    LocalMux I__10264 (
            .O(N__45159),
            .I(N__45150));
    Sp12to4 I__10263 (
            .O(N__45156),
            .I(N__45147));
    Span4Mux_v I__10262 (
            .O(N__45153),
            .I(N__45144));
    Span4Mux_h I__10261 (
            .O(N__45150),
            .I(N__45141));
    Odrv12 I__10260 (
            .O(N__45147),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__10259 (
            .O(N__45144),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__10258 (
            .O(N__45141),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__10257 (
            .O(N__45134),
            .I(N__45131));
    LocalMux I__10256 (
            .O(N__45131),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__10255 (
            .O(N__45128),
            .I(N__45122));
    InMux I__10254 (
            .O(N__45127),
            .I(N__45122));
    LocalMux I__10253 (
            .O(N__45122),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    CEMux I__10252 (
            .O(N__45119),
            .I(N__45092));
    CEMux I__10251 (
            .O(N__45118),
            .I(N__45092));
    CEMux I__10250 (
            .O(N__45117),
            .I(N__45092));
    CEMux I__10249 (
            .O(N__45116),
            .I(N__45092));
    CEMux I__10248 (
            .O(N__45115),
            .I(N__45092));
    CEMux I__10247 (
            .O(N__45114),
            .I(N__45092));
    CEMux I__10246 (
            .O(N__45113),
            .I(N__45092));
    CEMux I__10245 (
            .O(N__45112),
            .I(N__45092));
    CEMux I__10244 (
            .O(N__45111),
            .I(N__45092));
    GlobalMux I__10243 (
            .O(N__45092),
            .I(N__45089));
    gio2CtrlBuf I__10242 (
            .O(N__45089),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    InMux I__10241 (
            .O(N__45086),
            .I(N__45082));
    CascadeMux I__10240 (
            .O(N__45085),
            .I(N__45078));
    LocalMux I__10239 (
            .O(N__45082),
            .I(N__45075));
    InMux I__10238 (
            .O(N__45081),
            .I(N__45072));
    InMux I__10237 (
            .O(N__45078),
            .I(N__45069));
    Span4Mux_h I__10236 (
            .O(N__45075),
            .I(N__45062));
    LocalMux I__10235 (
            .O(N__45072),
            .I(N__45062));
    LocalMux I__10234 (
            .O(N__45069),
            .I(N__45062));
    Odrv4 I__10233 (
            .O(N__45062),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    CascadeMux I__10232 (
            .O(N__45059),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__10231 (
            .O(N__45056),
            .I(N__45052));
    CascadeMux I__10230 (
            .O(N__45055),
            .I(N__45049));
    LocalMux I__10229 (
            .O(N__45052),
            .I(N__45046));
    InMux I__10228 (
            .O(N__45049),
            .I(N__45043));
    Span4Mux_v I__10227 (
            .O(N__45046),
            .I(N__45038));
    LocalMux I__10226 (
            .O(N__45043),
            .I(N__45038));
    Odrv4 I__10225 (
            .O(N__45038),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__10224 (
            .O(N__45035),
            .I(N__45032));
    LocalMux I__10223 (
            .O(N__45032),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__10222 (
            .O(N__45029),
            .I(N__45025));
    CascadeMux I__10221 (
            .O(N__45028),
            .I(N__45020));
    LocalMux I__10220 (
            .O(N__45025),
            .I(N__45017));
    InMux I__10219 (
            .O(N__45024),
            .I(N__45012));
    InMux I__10218 (
            .O(N__45023),
            .I(N__45012));
    InMux I__10217 (
            .O(N__45020),
            .I(N__45009));
    Span4Mux_v I__10216 (
            .O(N__45017),
            .I(N__45004));
    LocalMux I__10215 (
            .O(N__45012),
            .I(N__45004));
    LocalMux I__10214 (
            .O(N__45009),
            .I(N__44998));
    Span4Mux_v I__10213 (
            .O(N__45004),
            .I(N__44998));
    InMux I__10212 (
            .O(N__45003),
            .I(N__44995));
    Odrv4 I__10211 (
            .O(N__44998),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__10210 (
            .O(N__44995),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__10209 (
            .O(N__44990),
            .I(N__44982));
    CascadeMux I__10208 (
            .O(N__44989),
            .I(N__44978));
    CascadeMux I__10207 (
            .O(N__44988),
            .I(N__44974));
    InMux I__10206 (
            .O(N__44987),
            .I(N__44953));
    InMux I__10205 (
            .O(N__44986),
            .I(N__44953));
    InMux I__10204 (
            .O(N__44985),
            .I(N__44938));
    InMux I__10203 (
            .O(N__44982),
            .I(N__44938));
    InMux I__10202 (
            .O(N__44981),
            .I(N__44938));
    InMux I__10201 (
            .O(N__44978),
            .I(N__44938));
    InMux I__10200 (
            .O(N__44977),
            .I(N__44938));
    InMux I__10199 (
            .O(N__44974),
            .I(N__44938));
    InMux I__10198 (
            .O(N__44973),
            .I(N__44938));
    CascadeMux I__10197 (
            .O(N__44972),
            .I(N__44931));
    CascadeMux I__10196 (
            .O(N__44971),
            .I(N__44927));
    CascadeMux I__10195 (
            .O(N__44970),
            .I(N__44923));
    CascadeMux I__10194 (
            .O(N__44969),
            .I(N__44919));
    CascadeMux I__10193 (
            .O(N__44968),
            .I(N__44914));
    CascadeMux I__10192 (
            .O(N__44967),
            .I(N__44910));
    CascadeMux I__10191 (
            .O(N__44966),
            .I(N__44906));
    InMux I__10190 (
            .O(N__44965),
            .I(N__44902));
    InMux I__10189 (
            .O(N__44964),
            .I(N__44895));
    InMux I__10188 (
            .O(N__44963),
            .I(N__44895));
    InMux I__10187 (
            .O(N__44962),
            .I(N__44895));
    InMux I__10186 (
            .O(N__44961),
            .I(N__44882));
    InMux I__10185 (
            .O(N__44960),
            .I(N__44882));
    InMux I__10184 (
            .O(N__44959),
            .I(N__44882));
    InMux I__10183 (
            .O(N__44958),
            .I(N__44882));
    LocalMux I__10182 (
            .O(N__44953),
            .I(N__44877));
    LocalMux I__10181 (
            .O(N__44938),
            .I(N__44877));
    InMux I__10180 (
            .O(N__44937),
            .I(N__44868));
    InMux I__10179 (
            .O(N__44936),
            .I(N__44868));
    InMux I__10178 (
            .O(N__44935),
            .I(N__44868));
    InMux I__10177 (
            .O(N__44934),
            .I(N__44868));
    InMux I__10176 (
            .O(N__44931),
            .I(N__44851));
    InMux I__10175 (
            .O(N__44930),
            .I(N__44851));
    InMux I__10174 (
            .O(N__44927),
            .I(N__44851));
    InMux I__10173 (
            .O(N__44926),
            .I(N__44851));
    InMux I__10172 (
            .O(N__44923),
            .I(N__44851));
    InMux I__10171 (
            .O(N__44922),
            .I(N__44851));
    InMux I__10170 (
            .O(N__44919),
            .I(N__44851));
    InMux I__10169 (
            .O(N__44918),
            .I(N__44851));
    InMux I__10168 (
            .O(N__44917),
            .I(N__44836));
    InMux I__10167 (
            .O(N__44914),
            .I(N__44836));
    InMux I__10166 (
            .O(N__44913),
            .I(N__44836));
    InMux I__10165 (
            .O(N__44910),
            .I(N__44836));
    InMux I__10164 (
            .O(N__44909),
            .I(N__44836));
    InMux I__10163 (
            .O(N__44906),
            .I(N__44836));
    InMux I__10162 (
            .O(N__44905),
            .I(N__44836));
    LocalMux I__10161 (
            .O(N__44902),
            .I(N__44826));
    LocalMux I__10160 (
            .O(N__44895),
            .I(N__44826));
    InMux I__10159 (
            .O(N__44894),
            .I(N__44817));
    InMux I__10158 (
            .O(N__44893),
            .I(N__44817));
    InMux I__10157 (
            .O(N__44892),
            .I(N__44817));
    InMux I__10156 (
            .O(N__44891),
            .I(N__44817));
    LocalMux I__10155 (
            .O(N__44882),
            .I(N__44810));
    Span4Mux_v I__10154 (
            .O(N__44877),
            .I(N__44801));
    LocalMux I__10153 (
            .O(N__44868),
            .I(N__44801));
    LocalMux I__10152 (
            .O(N__44851),
            .I(N__44801));
    LocalMux I__10151 (
            .O(N__44836),
            .I(N__44801));
    InMux I__10150 (
            .O(N__44835),
            .I(N__44798));
    InMux I__10149 (
            .O(N__44834),
            .I(N__44793));
    InMux I__10148 (
            .O(N__44833),
            .I(N__44793));
    InMux I__10147 (
            .O(N__44832),
            .I(N__44790));
    InMux I__10146 (
            .O(N__44831),
            .I(N__44787));
    Span4Mux_v I__10145 (
            .O(N__44826),
            .I(N__44782));
    LocalMux I__10144 (
            .O(N__44817),
            .I(N__44779));
    InMux I__10143 (
            .O(N__44816),
            .I(N__44776));
    InMux I__10142 (
            .O(N__44815),
            .I(N__44771));
    InMux I__10141 (
            .O(N__44814),
            .I(N__44771));
    InMux I__10140 (
            .O(N__44813),
            .I(N__44768));
    Span4Mux_v I__10139 (
            .O(N__44810),
            .I(N__44763));
    Span4Mux_v I__10138 (
            .O(N__44801),
            .I(N__44763));
    LocalMux I__10137 (
            .O(N__44798),
            .I(N__44754));
    LocalMux I__10136 (
            .O(N__44793),
            .I(N__44754));
    LocalMux I__10135 (
            .O(N__44790),
            .I(N__44754));
    LocalMux I__10134 (
            .O(N__44787),
            .I(N__44754));
    InMux I__10133 (
            .O(N__44786),
            .I(N__44751));
    InMux I__10132 (
            .O(N__44785),
            .I(N__44748));
    Span4Mux_h I__10131 (
            .O(N__44782),
            .I(N__44735));
    Span4Mux_v I__10130 (
            .O(N__44779),
            .I(N__44735));
    LocalMux I__10129 (
            .O(N__44776),
            .I(N__44735));
    LocalMux I__10128 (
            .O(N__44771),
            .I(N__44735));
    LocalMux I__10127 (
            .O(N__44768),
            .I(N__44735));
    Sp12to4 I__10126 (
            .O(N__44763),
            .I(N__44730));
    Span12Mux_s11_v I__10125 (
            .O(N__44754),
            .I(N__44730));
    LocalMux I__10124 (
            .O(N__44751),
            .I(N__44727));
    LocalMux I__10123 (
            .O(N__44748),
            .I(N__44724));
    InMux I__10122 (
            .O(N__44747),
            .I(N__44721));
    CascadeMux I__10121 (
            .O(N__44746),
            .I(N__44717));
    Sp12to4 I__10120 (
            .O(N__44735),
            .I(N__44705));
    Span12Mux_h I__10119 (
            .O(N__44730),
            .I(N__44702));
    Span4Mux_s1_h I__10118 (
            .O(N__44727),
            .I(N__44695));
    Span4Mux_s1_v I__10117 (
            .O(N__44724),
            .I(N__44695));
    LocalMux I__10116 (
            .O(N__44721),
            .I(N__44695));
    InMux I__10115 (
            .O(N__44720),
            .I(N__44688));
    InMux I__10114 (
            .O(N__44717),
            .I(N__44688));
    InMux I__10113 (
            .O(N__44716),
            .I(N__44688));
    InMux I__10112 (
            .O(N__44715),
            .I(N__44685));
    InMux I__10111 (
            .O(N__44714),
            .I(N__44678));
    InMux I__10110 (
            .O(N__44713),
            .I(N__44678));
    InMux I__10109 (
            .O(N__44712),
            .I(N__44678));
    InMux I__10108 (
            .O(N__44711),
            .I(N__44669));
    InMux I__10107 (
            .O(N__44710),
            .I(N__44669));
    InMux I__10106 (
            .O(N__44709),
            .I(N__44669));
    InMux I__10105 (
            .O(N__44708),
            .I(N__44669));
    Span12Mux_v I__10104 (
            .O(N__44705),
            .I(N__44660));
    Span12Mux_h I__10103 (
            .O(N__44702),
            .I(N__44660));
    Sp12to4 I__10102 (
            .O(N__44695),
            .I(N__44660));
    LocalMux I__10101 (
            .O(N__44688),
            .I(N__44660));
    LocalMux I__10100 (
            .O(N__44685),
            .I(CONSTANT_ONE_NET));
    LocalMux I__10099 (
            .O(N__44678),
            .I(CONSTANT_ONE_NET));
    LocalMux I__10098 (
            .O(N__44669),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__10097 (
            .O(N__44660),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__10096 (
            .O(N__44651),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    CascadeMux I__10095 (
            .O(N__44648),
            .I(N__44645));
    InMux I__10094 (
            .O(N__44645),
            .I(N__44642));
    LocalMux I__10093 (
            .O(N__44642),
            .I(N__44638));
    InMux I__10092 (
            .O(N__44641),
            .I(N__44635));
    Span4Mux_h I__10091 (
            .O(N__44638),
            .I(N__44632));
    LocalMux I__10090 (
            .O(N__44635),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__10089 (
            .O(N__44632),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__10088 (
            .O(N__44627),
            .I(N__44624));
    LocalMux I__10087 (
            .O(N__44624),
            .I(N__44620));
    InMux I__10086 (
            .O(N__44623),
            .I(N__44617));
    Span4Mux_v I__10085 (
            .O(N__44620),
            .I(N__44612));
    LocalMux I__10084 (
            .O(N__44617),
            .I(N__44612));
    Span4Mux_h I__10083 (
            .O(N__44612),
            .I(N__44609));
    Odrv4 I__10082 (
            .O(N__44609),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__10081 (
            .O(N__44606),
            .I(N__44602));
    InMux I__10080 (
            .O(N__44605),
            .I(N__44599));
    LocalMux I__10079 (
            .O(N__44602),
            .I(N__44595));
    LocalMux I__10078 (
            .O(N__44599),
            .I(N__44592));
    InMux I__10077 (
            .O(N__44598),
            .I(N__44589));
    Span4Mux_h I__10076 (
            .O(N__44595),
            .I(N__44586));
    Odrv12 I__10075 (
            .O(N__44592),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__10074 (
            .O(N__44589),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__10073 (
            .O(N__44586),
            .I(\current_shift_inst.un4_control_input1_12 ));
    CascadeMux I__10072 (
            .O(N__44579),
            .I(N__44576));
    InMux I__10071 (
            .O(N__44576),
            .I(N__44573));
    LocalMux I__10070 (
            .O(N__44573),
            .I(N__44570));
    Span4Mux_h I__10069 (
            .O(N__44570),
            .I(N__44567));
    Odrv4 I__10068 (
            .O(N__44567),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__10067 (
            .O(N__44564),
            .I(N__44561));
    LocalMux I__10066 (
            .O(N__44561),
            .I(N__44558));
    Span4Mux_v I__10065 (
            .O(N__44558),
            .I(N__44555));
    Odrv4 I__10064 (
            .O(N__44555),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__10063 (
            .O(N__44552),
            .I(N__44548));
    InMux I__10062 (
            .O(N__44551),
            .I(N__44545));
    LocalMux I__10061 (
            .O(N__44548),
            .I(N__44542));
    LocalMux I__10060 (
            .O(N__44545),
            .I(N__44538));
    Span4Mux_h I__10059 (
            .O(N__44542),
            .I(N__44535));
    InMux I__10058 (
            .O(N__44541),
            .I(N__44532));
    Odrv12 I__10057 (
            .O(N__44538),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv4 I__10056 (
            .O(N__44535),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__10055 (
            .O(N__44532),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__10054 (
            .O(N__44525),
            .I(N__44522));
    LocalMux I__10053 (
            .O(N__44522),
            .I(N__44519));
    Odrv12 I__10052 (
            .O(N__44519),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ));
    InMux I__10051 (
            .O(N__44516),
            .I(N__44513));
    LocalMux I__10050 (
            .O(N__44513),
            .I(N__44509));
    InMux I__10049 (
            .O(N__44512),
            .I(N__44506));
    Span4Mux_v I__10048 (
            .O(N__44509),
            .I(N__44500));
    LocalMux I__10047 (
            .O(N__44506),
            .I(N__44500));
    InMux I__10046 (
            .O(N__44505),
            .I(N__44496));
    Span4Mux_v I__10045 (
            .O(N__44500),
            .I(N__44493));
    InMux I__10044 (
            .O(N__44499),
            .I(N__44490));
    LocalMux I__10043 (
            .O(N__44496),
            .I(N__44487));
    Odrv4 I__10042 (
            .O(N__44493),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__10041 (
            .O(N__44490),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__10040 (
            .O(N__44487),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__10039 (
            .O(N__44480),
            .I(N__44477));
    LocalMux I__10038 (
            .O(N__44477),
            .I(N__44474));
    Span4Mux_v I__10037 (
            .O(N__44474),
            .I(N__44470));
    InMux I__10036 (
            .O(N__44473),
            .I(N__44467));
    Span4Mux_v I__10035 (
            .O(N__44470),
            .I(N__44461));
    LocalMux I__10034 (
            .O(N__44467),
            .I(N__44461));
    InMux I__10033 (
            .O(N__44466),
            .I(N__44458));
    Span4Mux_h I__10032 (
            .O(N__44461),
            .I(N__44455));
    LocalMux I__10031 (
            .O(N__44458),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__10030 (
            .O(N__44455),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    CascadeMux I__10029 (
            .O(N__44450),
            .I(N__44447));
    InMux I__10028 (
            .O(N__44447),
            .I(N__44444));
    LocalMux I__10027 (
            .O(N__44444),
            .I(N__44441));
    Odrv12 I__10026 (
            .O(N__44441),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    InMux I__10025 (
            .O(N__44438),
            .I(N__44431));
    InMux I__10024 (
            .O(N__44437),
            .I(N__44431));
    InMux I__10023 (
            .O(N__44436),
            .I(N__44428));
    LocalMux I__10022 (
            .O(N__44431),
            .I(N__44425));
    LocalMux I__10021 (
            .O(N__44428),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv12 I__10020 (
            .O(N__44425),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    CascadeMux I__10019 (
            .O(N__44420),
            .I(N__44417));
    InMux I__10018 (
            .O(N__44417),
            .I(N__44411));
    InMux I__10017 (
            .O(N__44416),
            .I(N__44411));
    LocalMux I__10016 (
            .O(N__44411),
            .I(N__44407));
    InMux I__10015 (
            .O(N__44410),
            .I(N__44404));
    Span4Mux_v I__10014 (
            .O(N__44407),
            .I(N__44401));
    LocalMux I__10013 (
            .O(N__44404),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__10012 (
            .O(N__44401),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__10011 (
            .O(N__44396),
            .I(N__44393));
    LocalMux I__10010 (
            .O(N__44393),
            .I(N__44390));
    Odrv12 I__10009 (
            .O(N__44390),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    InMux I__10008 (
            .O(N__44387),
            .I(N__44382));
    InMux I__10007 (
            .O(N__44386),
            .I(N__44379));
    InMux I__10006 (
            .O(N__44385),
            .I(N__44376));
    LocalMux I__10005 (
            .O(N__44382),
            .I(N__44371));
    LocalMux I__10004 (
            .O(N__44379),
            .I(N__44371));
    LocalMux I__10003 (
            .O(N__44376),
            .I(N__44368));
    Span4Mux_v I__10002 (
            .O(N__44371),
            .I(N__44365));
    Span4Mux_v I__10001 (
            .O(N__44368),
            .I(N__44359));
    Span4Mux_h I__10000 (
            .O(N__44365),
            .I(N__44359));
    InMux I__9999 (
            .O(N__44364),
            .I(N__44356));
    Odrv4 I__9998 (
            .O(N__44359),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__9997 (
            .O(N__44356),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__9996 (
            .O(N__44351),
            .I(N__44348));
    LocalMux I__9995 (
            .O(N__44348),
            .I(N__44345));
    Span4Mux_v I__9994 (
            .O(N__44345),
            .I(N__44342));
    Span4Mux_h I__9993 (
            .O(N__44342),
            .I(N__44337));
    InMux I__9992 (
            .O(N__44341),
            .I(N__44334));
    InMux I__9991 (
            .O(N__44340),
            .I(N__44331));
    Span4Mux_h I__9990 (
            .O(N__44337),
            .I(N__44328));
    LocalMux I__9989 (
            .O(N__44334),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    LocalMux I__9988 (
            .O(N__44331),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    Odrv4 I__9987 (
            .O(N__44328),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__9986 (
            .O(N__44321),
            .I(N__44315));
    InMux I__9985 (
            .O(N__44320),
            .I(N__44315));
    LocalMux I__9984 (
            .O(N__44315),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    InMux I__9983 (
            .O(N__44312),
            .I(N__44309));
    LocalMux I__9982 (
            .O(N__44309),
            .I(N__44306));
    Span4Mux_h I__9981 (
            .O(N__44306),
            .I(N__44302));
    InMux I__9980 (
            .O(N__44305),
            .I(N__44299));
    Span4Mux_v I__9979 (
            .O(N__44302),
            .I(N__44295));
    LocalMux I__9978 (
            .O(N__44299),
            .I(N__44292));
    InMux I__9977 (
            .O(N__44298),
            .I(N__44289));
    Span4Mux_h I__9976 (
            .O(N__44295),
            .I(N__44286));
    Span4Mux_s2_v I__9975 (
            .O(N__44292),
            .I(N__44283));
    LocalMux I__9974 (
            .O(N__44289),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__9973 (
            .O(N__44286),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__9972 (
            .O(N__44283),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__9971 (
            .O(N__44276),
            .I(N__44273));
    LocalMux I__9970 (
            .O(N__44273),
            .I(N__44268));
    InMux I__9969 (
            .O(N__44272),
            .I(N__44265));
    InMux I__9968 (
            .O(N__44271),
            .I(N__44262));
    Span4Mux_v I__9967 (
            .O(N__44268),
            .I(N__44257));
    LocalMux I__9966 (
            .O(N__44265),
            .I(N__44257));
    LocalMux I__9965 (
            .O(N__44262),
            .I(N__44253));
    Span4Mux_v I__9964 (
            .O(N__44257),
            .I(N__44250));
    CascadeMux I__9963 (
            .O(N__44256),
            .I(N__44247));
    Span4Mux_v I__9962 (
            .O(N__44253),
            .I(N__44244));
    Span4Mux_h I__9961 (
            .O(N__44250),
            .I(N__44241));
    InMux I__9960 (
            .O(N__44247),
            .I(N__44238));
    Odrv4 I__9959 (
            .O(N__44244),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__9958 (
            .O(N__44241),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__9957 (
            .O(N__44238),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    CascadeMux I__9956 (
            .O(N__44231),
            .I(N__44228));
    InMux I__9955 (
            .O(N__44228),
            .I(N__44222));
    InMux I__9954 (
            .O(N__44227),
            .I(N__44222));
    LocalMux I__9953 (
            .O(N__44222),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    InMux I__9952 (
            .O(N__44219),
            .I(N__44216));
    LocalMux I__9951 (
            .O(N__44216),
            .I(N__44213));
    Odrv4 I__9950 (
            .O(N__44213),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    InMux I__9949 (
            .O(N__44210),
            .I(N__44204));
    InMux I__9948 (
            .O(N__44209),
            .I(N__44204));
    LocalMux I__9947 (
            .O(N__44204),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    CascadeMux I__9946 (
            .O(N__44201),
            .I(N__44197));
    InMux I__9945 (
            .O(N__44200),
            .I(N__44192));
    InMux I__9944 (
            .O(N__44197),
            .I(N__44192));
    LocalMux I__9943 (
            .O(N__44192),
            .I(N__44188));
    InMux I__9942 (
            .O(N__44191),
            .I(N__44185));
    Span4Mux_v I__9941 (
            .O(N__44188),
            .I(N__44182));
    LocalMux I__9940 (
            .O(N__44185),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__9939 (
            .O(N__44182),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    CascadeMux I__9938 (
            .O(N__44177),
            .I(N__44173));
    InMux I__9937 (
            .O(N__44176),
            .I(N__44168));
    InMux I__9936 (
            .O(N__44173),
            .I(N__44168));
    LocalMux I__9935 (
            .O(N__44168),
            .I(N__44164));
    InMux I__9934 (
            .O(N__44167),
            .I(N__44161));
    Span4Mux_h I__9933 (
            .O(N__44164),
            .I(N__44158));
    LocalMux I__9932 (
            .O(N__44161),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__9931 (
            .O(N__44158),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__9930 (
            .O(N__44153),
            .I(N__44150));
    InMux I__9929 (
            .O(N__44150),
            .I(N__44147));
    LocalMux I__9928 (
            .O(N__44147),
            .I(N__44144));
    Odrv12 I__9927 (
            .O(N__44144),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    InMux I__9926 (
            .O(N__44141),
            .I(N__44133));
    InMux I__9925 (
            .O(N__44140),
            .I(N__44133));
    InMux I__9924 (
            .O(N__44139),
            .I(N__44130));
    InMux I__9923 (
            .O(N__44138),
            .I(N__44127));
    LocalMux I__9922 (
            .O(N__44133),
            .I(N__44122));
    LocalMux I__9921 (
            .O(N__44130),
            .I(N__44122));
    LocalMux I__9920 (
            .O(N__44127),
            .I(N__44119));
    Span4Mux_v I__9919 (
            .O(N__44122),
            .I(N__44116));
    Odrv12 I__9918 (
            .O(N__44119),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__9917 (
            .O(N__44116),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__9916 (
            .O(N__44111),
            .I(N__44108));
    LocalMux I__9915 (
            .O(N__44108),
            .I(N__44105));
    Span4Mux_v I__9914 (
            .O(N__44105),
            .I(N__44102));
    Span4Mux_v I__9913 (
            .O(N__44102),
            .I(N__44098));
    InMux I__9912 (
            .O(N__44101),
            .I(N__44095));
    Odrv4 I__9911 (
            .O(N__44098),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    LocalMux I__9910 (
            .O(N__44095),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    CascadeMux I__9909 (
            .O(N__44090),
            .I(N__44087));
    InMux I__9908 (
            .O(N__44087),
            .I(N__44083));
    InMux I__9907 (
            .O(N__44086),
            .I(N__44080));
    LocalMux I__9906 (
            .O(N__44083),
            .I(N__44074));
    LocalMux I__9905 (
            .O(N__44080),
            .I(N__44074));
    InMux I__9904 (
            .O(N__44079),
            .I(N__44071));
    Span4Mux_h I__9903 (
            .O(N__44074),
            .I(N__44068));
    LocalMux I__9902 (
            .O(N__44071),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__9901 (
            .O(N__44068),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__9900 (
            .O(N__44063),
            .I(N__44060));
    LocalMux I__9899 (
            .O(N__44060),
            .I(N__44055));
    InMux I__9898 (
            .O(N__44059),
            .I(N__44052));
    InMux I__9897 (
            .O(N__44058),
            .I(N__44049));
    Span4Mux_v I__9896 (
            .O(N__44055),
            .I(N__44044));
    LocalMux I__9895 (
            .O(N__44052),
            .I(N__44044));
    LocalMux I__9894 (
            .O(N__44049),
            .I(N__44041));
    Span4Mux_h I__9893 (
            .O(N__44044),
            .I(N__44038));
    Span4Mux_h I__9892 (
            .O(N__44041),
            .I(N__44034));
    Span4Mux_v I__9891 (
            .O(N__44038),
            .I(N__44031));
    InMux I__9890 (
            .O(N__44037),
            .I(N__44028));
    Odrv4 I__9889 (
            .O(N__44034),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__9888 (
            .O(N__44031),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__9887 (
            .O(N__44028),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__9886 (
            .O(N__44021),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__9885 (
            .O(N__44018),
            .I(N__44015));
    InMux I__9884 (
            .O(N__44015),
            .I(N__44011));
    InMux I__9883 (
            .O(N__44014),
            .I(N__44008));
    LocalMux I__9882 (
            .O(N__44011),
            .I(N__44004));
    LocalMux I__9881 (
            .O(N__44008),
            .I(N__44001));
    InMux I__9880 (
            .O(N__44007),
            .I(N__43998));
    Span4Mux_h I__9879 (
            .O(N__44004),
            .I(N__43995));
    Span4Mux_h I__9878 (
            .O(N__44001),
            .I(N__43992));
    LocalMux I__9877 (
            .O(N__43998),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__9876 (
            .O(N__43995),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__9875 (
            .O(N__43992),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__9874 (
            .O(N__43985),
            .I(N__43980));
    InMux I__9873 (
            .O(N__43984),
            .I(N__43977));
    InMux I__9872 (
            .O(N__43983),
            .I(N__43974));
    LocalMux I__9871 (
            .O(N__43980),
            .I(N__43969));
    LocalMux I__9870 (
            .O(N__43977),
            .I(N__43969));
    LocalMux I__9869 (
            .O(N__43974),
            .I(N__43965));
    Span4Mux_v I__9868 (
            .O(N__43969),
            .I(N__43962));
    InMux I__9867 (
            .O(N__43968),
            .I(N__43959));
    Span4Mux_v I__9866 (
            .O(N__43965),
            .I(N__43956));
    Span4Mux_h I__9865 (
            .O(N__43962),
            .I(N__43951));
    LocalMux I__9864 (
            .O(N__43959),
            .I(N__43951));
    Odrv4 I__9863 (
            .O(N__43956),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__9862 (
            .O(N__43951),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__9861 (
            .O(N__43946),
            .I(bfn_18_10_0_));
    CascadeMux I__9860 (
            .O(N__43943),
            .I(N__43939));
    InMux I__9859 (
            .O(N__43942),
            .I(N__43936));
    InMux I__9858 (
            .O(N__43939),
            .I(N__43932));
    LocalMux I__9857 (
            .O(N__43936),
            .I(N__43929));
    InMux I__9856 (
            .O(N__43935),
            .I(N__43926));
    LocalMux I__9855 (
            .O(N__43932),
            .I(N__43923));
    Span4Mux_h I__9854 (
            .O(N__43929),
            .I(N__43920));
    LocalMux I__9853 (
            .O(N__43926),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__9852 (
            .O(N__43923),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__9851 (
            .O(N__43920),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__9850 (
            .O(N__43913),
            .I(N__43906));
    InMux I__9849 (
            .O(N__43912),
            .I(N__43906));
    InMux I__9848 (
            .O(N__43911),
            .I(N__43902));
    LocalMux I__9847 (
            .O(N__43906),
            .I(N__43899));
    InMux I__9846 (
            .O(N__43905),
            .I(N__43896));
    LocalMux I__9845 (
            .O(N__43902),
            .I(N__43893));
    Span4Mux_h I__9844 (
            .O(N__43899),
            .I(N__43890));
    LocalMux I__9843 (
            .O(N__43896),
            .I(N__43887));
    Odrv4 I__9842 (
            .O(N__43893),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__9841 (
            .O(N__43890),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__9840 (
            .O(N__43887),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__9839 (
            .O(N__43880),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__9838 (
            .O(N__43877),
            .I(N__43870));
    InMux I__9837 (
            .O(N__43876),
            .I(N__43870));
    InMux I__9836 (
            .O(N__43875),
            .I(N__43867));
    LocalMux I__9835 (
            .O(N__43870),
            .I(N__43864));
    LocalMux I__9834 (
            .O(N__43867),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv4 I__9833 (
            .O(N__43864),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    CascadeMux I__9832 (
            .O(N__43859),
            .I(N__43856));
    InMux I__9831 (
            .O(N__43856),
            .I(N__43852));
    InMux I__9830 (
            .O(N__43855),
            .I(N__43849));
    LocalMux I__9829 (
            .O(N__43852),
            .I(N__43846));
    LocalMux I__9828 (
            .O(N__43849),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__9827 (
            .O(N__43846),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__9826 (
            .O(N__43841),
            .I(N__43834));
    InMux I__9825 (
            .O(N__43840),
            .I(N__43834));
    InMux I__9824 (
            .O(N__43839),
            .I(N__43831));
    LocalMux I__9823 (
            .O(N__43834),
            .I(N__43828));
    LocalMux I__9822 (
            .O(N__43831),
            .I(N__43824));
    Span4Mux_h I__9821 (
            .O(N__43828),
            .I(N__43821));
    InMux I__9820 (
            .O(N__43827),
            .I(N__43818));
    Odrv4 I__9819 (
            .O(N__43824),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    Odrv4 I__9818 (
            .O(N__43821),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__9817 (
            .O(N__43818),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__9816 (
            .O(N__43811),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__9815 (
            .O(N__43808),
            .I(N__43805));
    LocalMux I__9814 (
            .O(N__43805),
            .I(N__43801));
    InMux I__9813 (
            .O(N__43804),
            .I(N__43798));
    Span4Mux_v I__9812 (
            .O(N__43801),
            .I(N__43795));
    LocalMux I__9811 (
            .O(N__43798),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__9810 (
            .O(N__43795),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__9809 (
            .O(N__43790),
            .I(N__43787));
    InMux I__9808 (
            .O(N__43787),
            .I(N__43783));
    InMux I__9807 (
            .O(N__43786),
            .I(N__43780));
    LocalMux I__9806 (
            .O(N__43783),
            .I(N__43774));
    LocalMux I__9805 (
            .O(N__43780),
            .I(N__43774));
    InMux I__9804 (
            .O(N__43779),
            .I(N__43771));
    Span4Mux_h I__9803 (
            .O(N__43774),
            .I(N__43768));
    LocalMux I__9802 (
            .O(N__43771),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv4 I__9801 (
            .O(N__43768),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__9800 (
            .O(N__43763),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__9799 (
            .O(N__43760),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__9798 (
            .O(N__43757),
            .I(N__43754));
    InMux I__9797 (
            .O(N__43754),
            .I(N__43751));
    LocalMux I__9796 (
            .O(N__43751),
            .I(N__43746));
    InMux I__9795 (
            .O(N__43750),
            .I(N__43743));
    InMux I__9794 (
            .O(N__43749),
            .I(N__43740));
    Span4Mux_h I__9793 (
            .O(N__43746),
            .I(N__43737));
    LocalMux I__9792 (
            .O(N__43743),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__9791 (
            .O(N__43740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__9790 (
            .O(N__43737),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    CascadeMux I__9789 (
            .O(N__43730),
            .I(N__43727));
    InMux I__9788 (
            .O(N__43727),
            .I(N__43724));
    LocalMux I__9787 (
            .O(N__43724),
            .I(N__43719));
    InMux I__9786 (
            .O(N__43723),
            .I(N__43716));
    InMux I__9785 (
            .O(N__43722),
            .I(N__43713));
    Span12Mux_s8_h I__9784 (
            .O(N__43719),
            .I(N__43710));
    LocalMux I__9783 (
            .O(N__43716),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__9782 (
            .O(N__43713),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv12 I__9781 (
            .O(N__43710),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__9780 (
            .O(N__43703),
            .I(N__43697));
    InMux I__9779 (
            .O(N__43702),
            .I(N__43694));
    InMux I__9778 (
            .O(N__43701),
            .I(N__43691));
    CascadeMux I__9777 (
            .O(N__43700),
            .I(N__43688));
    LocalMux I__9776 (
            .O(N__43697),
            .I(N__43685));
    LocalMux I__9775 (
            .O(N__43694),
            .I(N__43682));
    LocalMux I__9774 (
            .O(N__43691),
            .I(N__43679));
    InMux I__9773 (
            .O(N__43688),
            .I(N__43676));
    Span4Mux_h I__9772 (
            .O(N__43685),
            .I(N__43671));
    Span4Mux_h I__9771 (
            .O(N__43682),
            .I(N__43671));
    Span4Mux_h I__9770 (
            .O(N__43679),
            .I(N__43668));
    LocalMux I__9769 (
            .O(N__43676),
            .I(N__43665));
    Sp12to4 I__9768 (
            .O(N__43671),
            .I(N__43662));
    Span4Mux_v I__9767 (
            .O(N__43668),
            .I(N__43657));
    Span4Mux_h I__9766 (
            .O(N__43665),
            .I(N__43657));
    Odrv12 I__9765 (
            .O(N__43662),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    Odrv4 I__9764 (
            .O(N__43657),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    CEMux I__9763 (
            .O(N__43652),
            .I(N__43646));
    CEMux I__9762 (
            .O(N__43651),
            .I(N__43642));
    CEMux I__9761 (
            .O(N__43650),
            .I(N__43639));
    CEMux I__9760 (
            .O(N__43649),
            .I(N__43636));
    LocalMux I__9759 (
            .O(N__43646),
            .I(N__43633));
    CEMux I__9758 (
            .O(N__43645),
            .I(N__43630));
    LocalMux I__9757 (
            .O(N__43642),
            .I(N__43627));
    LocalMux I__9756 (
            .O(N__43639),
            .I(N__43624));
    LocalMux I__9755 (
            .O(N__43636),
            .I(N__43621));
    Span4Mux_h I__9754 (
            .O(N__43633),
            .I(N__43618));
    LocalMux I__9753 (
            .O(N__43630),
            .I(N__43615));
    Span4Mux_v I__9752 (
            .O(N__43627),
            .I(N__43612));
    Span4Mux_v I__9751 (
            .O(N__43624),
            .I(N__43609));
    Span4Mux_v I__9750 (
            .O(N__43621),
            .I(N__43606));
    Span4Mux_h I__9749 (
            .O(N__43618),
            .I(N__43603));
    Span4Mux_h I__9748 (
            .O(N__43615),
            .I(N__43600));
    Span4Mux_h I__9747 (
            .O(N__43612),
            .I(N__43595));
    Span4Mux_h I__9746 (
            .O(N__43609),
            .I(N__43595));
    Span4Mux_h I__9745 (
            .O(N__43606),
            .I(N__43592));
    Span4Mux_v I__9744 (
            .O(N__43603),
            .I(N__43587));
    Span4Mux_h I__9743 (
            .O(N__43600),
            .I(N__43587));
    Odrv4 I__9742 (
            .O(N__43595),
            .I(\delay_measurement_inst.delay_hc_timer.N_163_i ));
    Odrv4 I__9741 (
            .O(N__43592),
            .I(\delay_measurement_inst.delay_hc_timer.N_163_i ));
    Odrv4 I__9740 (
            .O(N__43587),
            .I(\delay_measurement_inst.delay_hc_timer.N_163_i ));
    InMux I__9739 (
            .O(N__43580),
            .I(N__43574));
    InMux I__9738 (
            .O(N__43579),
            .I(N__43574));
    LocalMux I__9737 (
            .O(N__43574),
            .I(N__43570));
    InMux I__9736 (
            .O(N__43573),
            .I(N__43567));
    Span4Mux_h I__9735 (
            .O(N__43570),
            .I(N__43564));
    LocalMux I__9734 (
            .O(N__43567),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__9733 (
            .O(N__43564),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__9732 (
            .O(N__43559),
            .I(N__43556));
    LocalMux I__9731 (
            .O(N__43556),
            .I(N__43551));
    InMux I__9730 (
            .O(N__43555),
            .I(N__43548));
    InMux I__9729 (
            .O(N__43554),
            .I(N__43545));
    Span4Mux_h I__9728 (
            .O(N__43551),
            .I(N__43541));
    LocalMux I__9727 (
            .O(N__43548),
            .I(N__43536));
    LocalMux I__9726 (
            .O(N__43545),
            .I(N__43536));
    InMux I__9725 (
            .O(N__43544),
            .I(N__43533));
    Odrv4 I__9724 (
            .O(N__43541),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv12 I__9723 (
            .O(N__43536),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__9722 (
            .O(N__43533),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__9721 (
            .O(N__43526),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__9720 (
            .O(N__43523),
            .I(N__43520));
    InMux I__9719 (
            .O(N__43520),
            .I(N__43516));
    InMux I__9718 (
            .O(N__43519),
            .I(N__43513));
    LocalMux I__9717 (
            .O(N__43516),
            .I(N__43509));
    LocalMux I__9716 (
            .O(N__43513),
            .I(N__43506));
    InMux I__9715 (
            .O(N__43512),
            .I(N__43503));
    Span4Mux_h I__9714 (
            .O(N__43509),
            .I(N__43500));
    Span4Mux_h I__9713 (
            .O(N__43506),
            .I(N__43497));
    LocalMux I__9712 (
            .O(N__43503),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__9711 (
            .O(N__43500),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__9710 (
            .O(N__43497),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__9709 (
            .O(N__43490),
            .I(N__43483));
    InMux I__9708 (
            .O(N__43489),
            .I(N__43483));
    InMux I__9707 (
            .O(N__43488),
            .I(N__43480));
    LocalMux I__9706 (
            .O(N__43483),
            .I(N__43477));
    LocalMux I__9705 (
            .O(N__43480),
            .I(N__43471));
    Span12Mux_s8_v I__9704 (
            .O(N__43477),
            .I(N__43471));
    InMux I__9703 (
            .O(N__43476),
            .I(N__43468));
    Odrv12 I__9702 (
            .O(N__43471),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    LocalMux I__9701 (
            .O(N__43468),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__9700 (
            .O(N__43463),
            .I(bfn_18_9_0_));
    CascadeMux I__9699 (
            .O(N__43460),
            .I(N__43456));
    CascadeMux I__9698 (
            .O(N__43459),
            .I(N__43453));
    InMux I__9697 (
            .O(N__43456),
            .I(N__43450));
    InMux I__9696 (
            .O(N__43453),
            .I(N__43446));
    LocalMux I__9695 (
            .O(N__43450),
            .I(N__43443));
    InMux I__9694 (
            .O(N__43449),
            .I(N__43440));
    LocalMux I__9693 (
            .O(N__43446),
            .I(N__43437));
    Span4Mux_h I__9692 (
            .O(N__43443),
            .I(N__43434));
    LocalMux I__9691 (
            .O(N__43440),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__9690 (
            .O(N__43437),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__9689 (
            .O(N__43434),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__9688 (
            .O(N__43427),
            .I(N__43422));
    InMux I__9687 (
            .O(N__43426),
            .I(N__43417));
    InMux I__9686 (
            .O(N__43425),
            .I(N__43417));
    LocalMux I__9685 (
            .O(N__43422),
            .I(N__43413));
    LocalMux I__9684 (
            .O(N__43417),
            .I(N__43410));
    CascadeMux I__9683 (
            .O(N__43416),
            .I(N__43407));
    Span4Mux_h I__9682 (
            .O(N__43413),
            .I(N__43404));
    Span12Mux_s8_v I__9681 (
            .O(N__43410),
            .I(N__43401));
    InMux I__9680 (
            .O(N__43407),
            .I(N__43398));
    Odrv4 I__9679 (
            .O(N__43404),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv12 I__9678 (
            .O(N__43401),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__9677 (
            .O(N__43398),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__9676 (
            .O(N__43391),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__9675 (
            .O(N__43388),
            .I(N__43381));
    InMux I__9674 (
            .O(N__43387),
            .I(N__43381));
    InMux I__9673 (
            .O(N__43386),
            .I(N__43378));
    LocalMux I__9672 (
            .O(N__43381),
            .I(N__43375));
    LocalMux I__9671 (
            .O(N__43378),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__9670 (
            .O(N__43375),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__9669 (
            .O(N__43370),
            .I(N__43365));
    InMux I__9668 (
            .O(N__43369),
            .I(N__43362));
    InMux I__9667 (
            .O(N__43368),
            .I(N__43359));
    LocalMux I__9666 (
            .O(N__43365),
            .I(N__43356));
    LocalMux I__9665 (
            .O(N__43362),
            .I(N__43351));
    LocalMux I__9664 (
            .O(N__43359),
            .I(N__43351));
    Span4Mux_v I__9663 (
            .O(N__43356),
            .I(N__43347));
    Span12Mux_s8_v I__9662 (
            .O(N__43351),
            .I(N__43344));
    InMux I__9661 (
            .O(N__43350),
            .I(N__43341));
    Odrv4 I__9660 (
            .O(N__43347),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv12 I__9659 (
            .O(N__43344),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__9658 (
            .O(N__43341),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__9657 (
            .O(N__43334),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__9656 (
            .O(N__43331),
            .I(N__43324));
    InMux I__9655 (
            .O(N__43330),
            .I(N__43324));
    InMux I__9654 (
            .O(N__43329),
            .I(N__43321));
    LocalMux I__9653 (
            .O(N__43324),
            .I(N__43318));
    LocalMux I__9652 (
            .O(N__43321),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv4 I__9651 (
            .O(N__43318),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__9650 (
            .O(N__43313),
            .I(N__43310));
    LocalMux I__9649 (
            .O(N__43310),
            .I(N__43305));
    InMux I__9648 (
            .O(N__43309),
            .I(N__43300));
    InMux I__9647 (
            .O(N__43308),
            .I(N__43300));
    Span4Mux_v I__9646 (
            .O(N__43305),
            .I(N__43294));
    LocalMux I__9645 (
            .O(N__43300),
            .I(N__43294));
    CascadeMux I__9644 (
            .O(N__43299),
            .I(N__43291));
    Span4Mux_v I__9643 (
            .O(N__43294),
            .I(N__43288));
    InMux I__9642 (
            .O(N__43291),
            .I(N__43285));
    Odrv4 I__9641 (
            .O(N__43288),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__9640 (
            .O(N__43285),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__9639 (
            .O(N__43280),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__9638 (
            .O(N__43277),
            .I(N__43273));
    CascadeMux I__9637 (
            .O(N__43276),
            .I(N__43270));
    InMux I__9636 (
            .O(N__43273),
            .I(N__43264));
    InMux I__9635 (
            .O(N__43270),
            .I(N__43264));
    InMux I__9634 (
            .O(N__43269),
            .I(N__43261));
    LocalMux I__9633 (
            .O(N__43264),
            .I(N__43258));
    LocalMux I__9632 (
            .O(N__43261),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__9631 (
            .O(N__43258),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__9630 (
            .O(N__43253),
            .I(N__43248));
    InMux I__9629 (
            .O(N__43252),
            .I(N__43243));
    InMux I__9628 (
            .O(N__43251),
            .I(N__43243));
    LocalMux I__9627 (
            .O(N__43248),
            .I(N__43240));
    LocalMux I__9626 (
            .O(N__43243),
            .I(N__43237));
    Span4Mux_h I__9625 (
            .O(N__43240),
            .I(N__43233));
    Span4Mux_h I__9624 (
            .O(N__43237),
            .I(N__43230));
    InMux I__9623 (
            .O(N__43236),
            .I(N__43227));
    Odrv4 I__9622 (
            .O(N__43233),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv4 I__9621 (
            .O(N__43230),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__9620 (
            .O(N__43227),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__9619 (
            .O(N__43220),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__9618 (
            .O(N__43217),
            .I(N__43213));
    CascadeMux I__9617 (
            .O(N__43216),
            .I(N__43210));
    InMux I__9616 (
            .O(N__43213),
            .I(N__43205));
    InMux I__9615 (
            .O(N__43210),
            .I(N__43205));
    LocalMux I__9614 (
            .O(N__43205),
            .I(N__43201));
    InMux I__9613 (
            .O(N__43204),
            .I(N__43198));
    Span4Mux_v I__9612 (
            .O(N__43201),
            .I(N__43195));
    LocalMux I__9611 (
            .O(N__43198),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__9610 (
            .O(N__43195),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__9609 (
            .O(N__43190),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__9608 (
            .O(N__43187),
            .I(N__43184));
    InMux I__9607 (
            .O(N__43184),
            .I(N__43180));
    InMux I__9606 (
            .O(N__43183),
            .I(N__43177));
    LocalMux I__9605 (
            .O(N__43180),
            .I(N__43171));
    LocalMux I__9604 (
            .O(N__43177),
            .I(N__43171));
    InMux I__9603 (
            .O(N__43176),
            .I(N__43168));
    Span4Mux_h I__9602 (
            .O(N__43171),
            .I(N__43165));
    LocalMux I__9601 (
            .O(N__43168),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__9600 (
            .O(N__43165),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__9599 (
            .O(N__43160),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__9598 (
            .O(N__43157),
            .I(N__43154));
    LocalMux I__9597 (
            .O(N__43154),
            .I(N__43151));
    Span4Mux_h I__9596 (
            .O(N__43151),
            .I(N__43147));
    CascadeMux I__9595 (
            .O(N__43150),
            .I(N__43142));
    Span4Mux_v I__9594 (
            .O(N__43147),
            .I(N__43139));
    InMux I__9593 (
            .O(N__43146),
            .I(N__43134));
    InMux I__9592 (
            .O(N__43145),
            .I(N__43134));
    InMux I__9591 (
            .O(N__43142),
            .I(N__43131));
    Odrv4 I__9590 (
            .O(N__43139),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__9589 (
            .O(N__43134),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__9588 (
            .O(N__43131),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__9587 (
            .O(N__43124),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__9586 (
            .O(N__43121),
            .I(N__43117));
    CascadeMux I__9585 (
            .O(N__43120),
            .I(N__43114));
    InMux I__9584 (
            .O(N__43117),
            .I(N__43111));
    InMux I__9583 (
            .O(N__43114),
            .I(N__43108));
    LocalMux I__9582 (
            .O(N__43111),
            .I(N__43104));
    LocalMux I__9581 (
            .O(N__43108),
            .I(N__43101));
    InMux I__9580 (
            .O(N__43107),
            .I(N__43098));
    Span4Mux_h I__9579 (
            .O(N__43104),
            .I(N__43095));
    Span4Mux_h I__9578 (
            .O(N__43101),
            .I(N__43092));
    LocalMux I__9577 (
            .O(N__43098),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__9576 (
            .O(N__43095),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__9575 (
            .O(N__43092),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__9574 (
            .O(N__43085),
            .I(N__43082));
    LocalMux I__9573 (
            .O(N__43082),
            .I(N__43079));
    Span4Mux_v I__9572 (
            .O(N__43079),
            .I(N__43073));
    InMux I__9571 (
            .O(N__43078),
            .I(N__43070));
    InMux I__9570 (
            .O(N__43077),
            .I(N__43065));
    InMux I__9569 (
            .O(N__43076),
            .I(N__43065));
    Odrv4 I__9568 (
            .O(N__43073),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__9567 (
            .O(N__43070),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__9566 (
            .O(N__43065),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__9565 (
            .O(N__43058),
            .I(bfn_18_8_0_));
    CascadeMux I__9564 (
            .O(N__43055),
            .I(N__43051));
    InMux I__9563 (
            .O(N__43054),
            .I(N__43048));
    InMux I__9562 (
            .O(N__43051),
            .I(N__43044));
    LocalMux I__9561 (
            .O(N__43048),
            .I(N__43041));
    InMux I__9560 (
            .O(N__43047),
            .I(N__43038));
    LocalMux I__9559 (
            .O(N__43044),
            .I(N__43033));
    Span4Mux_h I__9558 (
            .O(N__43041),
            .I(N__43033));
    LocalMux I__9557 (
            .O(N__43038),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__9556 (
            .O(N__43033),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__9555 (
            .O(N__43028),
            .I(N__43025));
    LocalMux I__9554 (
            .O(N__43025),
            .I(N__43021));
    InMux I__9553 (
            .O(N__43024),
            .I(N__43018));
    Span4Mux_v I__9552 (
            .O(N__43021),
            .I(N__43013));
    LocalMux I__9551 (
            .O(N__43018),
            .I(N__43010));
    InMux I__9550 (
            .O(N__43017),
            .I(N__43005));
    InMux I__9549 (
            .O(N__43016),
            .I(N__43005));
    Odrv4 I__9548 (
            .O(N__43013),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__9547 (
            .O(N__43010),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__9546 (
            .O(N__43005),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__9545 (
            .O(N__42998),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__9544 (
            .O(N__42995),
            .I(N__42988));
    InMux I__9543 (
            .O(N__42994),
            .I(N__42988));
    InMux I__9542 (
            .O(N__42993),
            .I(N__42985));
    LocalMux I__9541 (
            .O(N__42988),
            .I(N__42982));
    LocalMux I__9540 (
            .O(N__42985),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__9539 (
            .O(N__42982),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__9538 (
            .O(N__42977),
            .I(N__42974));
    LocalMux I__9537 (
            .O(N__42974),
            .I(N__42968));
    InMux I__9536 (
            .O(N__42973),
            .I(N__42963));
    InMux I__9535 (
            .O(N__42972),
            .I(N__42963));
    InMux I__9534 (
            .O(N__42971),
            .I(N__42960));
    Odrv4 I__9533 (
            .O(N__42968),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__9532 (
            .O(N__42963),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__9531 (
            .O(N__42960),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__9530 (
            .O(N__42953),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__9529 (
            .O(N__42950),
            .I(N__42943));
    InMux I__9528 (
            .O(N__42949),
            .I(N__42943));
    InMux I__9527 (
            .O(N__42948),
            .I(N__42940));
    LocalMux I__9526 (
            .O(N__42943),
            .I(N__42937));
    LocalMux I__9525 (
            .O(N__42940),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__9524 (
            .O(N__42937),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__9523 (
            .O(N__42932),
            .I(N__42929));
    LocalMux I__9522 (
            .O(N__42929),
            .I(N__42924));
    InMux I__9521 (
            .O(N__42928),
            .I(N__42921));
    InMux I__9520 (
            .O(N__42927),
            .I(N__42918));
    Span4Mux_h I__9519 (
            .O(N__42924),
            .I(N__42914));
    LocalMux I__9518 (
            .O(N__42921),
            .I(N__42909));
    LocalMux I__9517 (
            .O(N__42918),
            .I(N__42909));
    InMux I__9516 (
            .O(N__42917),
            .I(N__42906));
    Odrv4 I__9515 (
            .O(N__42914),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__9514 (
            .O(N__42909),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    LocalMux I__9513 (
            .O(N__42906),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__9512 (
            .O(N__42899),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__9511 (
            .O(N__42896),
            .I(N__42892));
    CascadeMux I__9510 (
            .O(N__42895),
            .I(N__42889));
    InMux I__9509 (
            .O(N__42892),
            .I(N__42883));
    InMux I__9508 (
            .O(N__42889),
            .I(N__42883));
    InMux I__9507 (
            .O(N__42888),
            .I(N__42880));
    LocalMux I__9506 (
            .O(N__42883),
            .I(N__42877));
    LocalMux I__9505 (
            .O(N__42880),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__9504 (
            .O(N__42877),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__9503 (
            .O(N__42872),
            .I(N__42869));
    LocalMux I__9502 (
            .O(N__42869),
            .I(N__42864));
    InMux I__9501 (
            .O(N__42868),
            .I(N__42859));
    InMux I__9500 (
            .O(N__42867),
            .I(N__42859));
    Span4Mux_v I__9499 (
            .O(N__42864),
            .I(N__42855));
    LocalMux I__9498 (
            .O(N__42859),
            .I(N__42852));
    InMux I__9497 (
            .O(N__42858),
            .I(N__42849));
    Odrv4 I__9496 (
            .O(N__42855),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv12 I__9495 (
            .O(N__42852),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    LocalMux I__9494 (
            .O(N__42849),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__9493 (
            .O(N__42842),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__9492 (
            .O(N__42839),
            .I(N__42835));
    CascadeMux I__9491 (
            .O(N__42838),
            .I(N__42832));
    InMux I__9490 (
            .O(N__42835),
            .I(N__42827));
    InMux I__9489 (
            .O(N__42832),
            .I(N__42827));
    LocalMux I__9488 (
            .O(N__42827),
            .I(N__42823));
    InMux I__9487 (
            .O(N__42826),
            .I(N__42820));
    Span4Mux_v I__9486 (
            .O(N__42823),
            .I(N__42817));
    LocalMux I__9485 (
            .O(N__42820),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__9484 (
            .O(N__42817),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__9483 (
            .O(N__42812),
            .I(N__42808));
    InMux I__9482 (
            .O(N__42811),
            .I(N__42805));
    LocalMux I__9481 (
            .O(N__42808),
            .I(N__42800));
    LocalMux I__9480 (
            .O(N__42805),
            .I(N__42797));
    InMux I__9479 (
            .O(N__42804),
            .I(N__42794));
    CascadeMux I__9478 (
            .O(N__42803),
            .I(N__42791));
    Span4Mux_v I__9477 (
            .O(N__42800),
            .I(N__42788));
    Span4Mux_h I__9476 (
            .O(N__42797),
            .I(N__42783));
    LocalMux I__9475 (
            .O(N__42794),
            .I(N__42783));
    InMux I__9474 (
            .O(N__42791),
            .I(N__42780));
    Odrv4 I__9473 (
            .O(N__42788),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__9472 (
            .O(N__42783),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__9471 (
            .O(N__42780),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__9470 (
            .O(N__42773),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__9469 (
            .O(N__42770),
            .I(N__42767));
    InMux I__9468 (
            .O(N__42767),
            .I(N__42763));
    InMux I__9467 (
            .O(N__42766),
            .I(N__42760));
    LocalMux I__9466 (
            .O(N__42763),
            .I(N__42754));
    LocalMux I__9465 (
            .O(N__42760),
            .I(N__42754));
    InMux I__9464 (
            .O(N__42759),
            .I(N__42751));
    Span4Mux_h I__9463 (
            .O(N__42754),
            .I(N__42748));
    LocalMux I__9462 (
            .O(N__42751),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__9461 (
            .O(N__42748),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__9460 (
            .O(N__42743),
            .I(N__42738));
    InMux I__9459 (
            .O(N__42742),
            .I(N__42733));
    InMux I__9458 (
            .O(N__42741),
            .I(N__42733));
    LocalMux I__9457 (
            .O(N__42738),
            .I(N__42730));
    LocalMux I__9456 (
            .O(N__42733),
            .I(N__42727));
    Span4Mux_h I__9455 (
            .O(N__42730),
            .I(N__42721));
    Span4Mux_h I__9454 (
            .O(N__42727),
            .I(N__42721));
    InMux I__9453 (
            .O(N__42726),
            .I(N__42718));
    Odrv4 I__9452 (
            .O(N__42721),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__9451 (
            .O(N__42718),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__9450 (
            .O(N__42713),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__9449 (
            .O(N__42710),
            .I(N__42706));
    InMux I__9448 (
            .O(N__42709),
            .I(N__42702));
    LocalMux I__9447 (
            .O(N__42706),
            .I(N__42699));
    InMux I__9446 (
            .O(N__42705),
            .I(N__42696));
    LocalMux I__9445 (
            .O(N__42702),
            .I(N__42691));
    Span4Mux_v I__9444 (
            .O(N__42699),
            .I(N__42691));
    LocalMux I__9443 (
            .O(N__42696),
            .I(N__42688));
    Odrv4 I__9442 (
            .O(N__42691),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv4 I__9441 (
            .O(N__42688),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    InMux I__9440 (
            .O(N__42683),
            .I(N__42680));
    LocalMux I__9439 (
            .O(N__42680),
            .I(N__42677));
    Span4Mux_h I__9438 (
            .O(N__42677),
            .I(N__42674));
    Odrv4 I__9437 (
            .O(N__42674),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__9436 (
            .O(N__42671),
            .I(N__42667));
    InMux I__9435 (
            .O(N__42670),
            .I(N__42663));
    LocalMux I__9434 (
            .O(N__42667),
            .I(N__42660));
    InMux I__9433 (
            .O(N__42666),
            .I(N__42657));
    LocalMux I__9432 (
            .O(N__42663),
            .I(N__42654));
    Span4Mux_h I__9431 (
            .O(N__42660),
            .I(N__42649));
    LocalMux I__9430 (
            .O(N__42657),
            .I(N__42649));
    Span4Mux_h I__9429 (
            .O(N__42654),
            .I(N__42643));
    Span4Mux_h I__9428 (
            .O(N__42649),
            .I(N__42643));
    InMux I__9427 (
            .O(N__42648),
            .I(N__42640));
    Odrv4 I__9426 (
            .O(N__42643),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__9425 (
            .O(N__42640),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__9424 (
            .O(N__42635),
            .I(N__42632));
    LocalMux I__9423 (
            .O(N__42632),
            .I(N__42627));
    InMux I__9422 (
            .O(N__42631),
            .I(N__42624));
    InMux I__9421 (
            .O(N__42630),
            .I(N__42621));
    Span4Mux_v I__9420 (
            .O(N__42627),
            .I(N__42618));
    LocalMux I__9419 (
            .O(N__42624),
            .I(N__42613));
    LocalMux I__9418 (
            .O(N__42621),
            .I(N__42613));
    Span4Mux_h I__9417 (
            .O(N__42618),
            .I(N__42607));
    Span4Mux_h I__9416 (
            .O(N__42613),
            .I(N__42607));
    InMux I__9415 (
            .O(N__42612),
            .I(N__42604));
    Odrv4 I__9414 (
            .O(N__42607),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__9413 (
            .O(N__42604),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__9412 (
            .O(N__42599),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__9411 (
            .O(N__42596),
            .I(N__42589));
    InMux I__9410 (
            .O(N__42595),
            .I(N__42589));
    InMux I__9409 (
            .O(N__42594),
            .I(N__42586));
    LocalMux I__9408 (
            .O(N__42589),
            .I(N__42583));
    LocalMux I__9407 (
            .O(N__42586),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__9406 (
            .O(N__42583),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__9405 (
            .O(N__42578),
            .I(N__42575));
    LocalMux I__9404 (
            .O(N__42575),
            .I(N__42570));
    InMux I__9403 (
            .O(N__42574),
            .I(N__42565));
    InMux I__9402 (
            .O(N__42573),
            .I(N__42565));
    Span4Mux_v I__9401 (
            .O(N__42570),
            .I(N__42560));
    LocalMux I__9400 (
            .O(N__42565),
            .I(N__42560));
    Span4Mux_h I__9399 (
            .O(N__42560),
            .I(N__42557));
    Span4Mux_h I__9398 (
            .O(N__42557),
            .I(N__42553));
    InMux I__9397 (
            .O(N__42556),
            .I(N__42550));
    Odrv4 I__9396 (
            .O(N__42553),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__9395 (
            .O(N__42550),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__9394 (
            .O(N__42545),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__9393 (
            .O(N__42542),
            .I(N__42535));
    InMux I__9392 (
            .O(N__42541),
            .I(N__42535));
    InMux I__9391 (
            .O(N__42540),
            .I(N__42532));
    LocalMux I__9390 (
            .O(N__42535),
            .I(N__42529));
    LocalMux I__9389 (
            .O(N__42532),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__9388 (
            .O(N__42529),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__9387 (
            .O(N__42524),
            .I(N__42521));
    LocalMux I__9386 (
            .O(N__42521),
            .I(N__42517));
    InMux I__9385 (
            .O(N__42520),
            .I(N__42514));
    Span4Mux_v I__9384 (
            .O(N__42517),
            .I(N__42510));
    LocalMux I__9383 (
            .O(N__42514),
            .I(N__42507));
    InMux I__9382 (
            .O(N__42513),
            .I(N__42504));
    Span4Mux_h I__9381 (
            .O(N__42510),
            .I(N__42500));
    Span4Mux_v I__9380 (
            .O(N__42507),
            .I(N__42497));
    LocalMux I__9379 (
            .O(N__42504),
            .I(N__42494));
    InMux I__9378 (
            .O(N__42503),
            .I(N__42491));
    Odrv4 I__9377 (
            .O(N__42500),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv4 I__9376 (
            .O(N__42497),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv12 I__9375 (
            .O(N__42494),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    LocalMux I__9374 (
            .O(N__42491),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__9373 (
            .O(N__42482),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__9372 (
            .O(N__42479),
            .I(N__42475));
    CascadeMux I__9371 (
            .O(N__42478),
            .I(N__42472));
    InMux I__9370 (
            .O(N__42475),
            .I(N__42466));
    InMux I__9369 (
            .O(N__42472),
            .I(N__42466));
    InMux I__9368 (
            .O(N__42471),
            .I(N__42463));
    LocalMux I__9367 (
            .O(N__42466),
            .I(N__42460));
    LocalMux I__9366 (
            .O(N__42463),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__9365 (
            .O(N__42460),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__9364 (
            .O(N__42455),
            .I(N__42451));
    InMux I__9363 (
            .O(N__42454),
            .I(N__42447));
    LocalMux I__9362 (
            .O(N__42451),
            .I(N__42444));
    InMux I__9361 (
            .O(N__42450),
            .I(N__42441));
    LocalMux I__9360 (
            .O(N__42447),
            .I(N__42438));
    Span4Mux_v I__9359 (
            .O(N__42444),
            .I(N__42433));
    LocalMux I__9358 (
            .O(N__42441),
            .I(N__42433));
    Span4Mux_v I__9357 (
            .O(N__42438),
            .I(N__42429));
    Span4Mux_h I__9356 (
            .O(N__42433),
            .I(N__42426));
    InMux I__9355 (
            .O(N__42432),
            .I(N__42423));
    Odrv4 I__9354 (
            .O(N__42429),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__9353 (
            .O(N__42426),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    LocalMux I__9352 (
            .O(N__42423),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__9351 (
            .O(N__42416),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__9350 (
            .O(N__42413),
            .I(N__42409));
    CascadeMux I__9349 (
            .O(N__42412),
            .I(N__42406));
    InMux I__9348 (
            .O(N__42409),
            .I(N__42400));
    InMux I__9347 (
            .O(N__42406),
            .I(N__42400));
    InMux I__9346 (
            .O(N__42405),
            .I(N__42397));
    LocalMux I__9345 (
            .O(N__42400),
            .I(N__42394));
    LocalMux I__9344 (
            .O(N__42397),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__9343 (
            .O(N__42394),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__9342 (
            .O(N__42389),
            .I(N__42385));
    InMux I__9341 (
            .O(N__42388),
            .I(N__42381));
    LocalMux I__9340 (
            .O(N__42385),
            .I(N__42378));
    InMux I__9339 (
            .O(N__42384),
            .I(N__42375));
    LocalMux I__9338 (
            .O(N__42381),
            .I(N__42372));
    Span4Mux_h I__9337 (
            .O(N__42378),
            .I(N__42369));
    LocalMux I__9336 (
            .O(N__42375),
            .I(N__42364));
    Span4Mux_h I__9335 (
            .O(N__42372),
            .I(N__42364));
    Span4Mux_h I__9334 (
            .O(N__42369),
            .I(N__42358));
    Span4Mux_h I__9333 (
            .O(N__42364),
            .I(N__42358));
    InMux I__9332 (
            .O(N__42363),
            .I(N__42355));
    Odrv4 I__9331 (
            .O(N__42358),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__9330 (
            .O(N__42355),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__9329 (
            .O(N__42350),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__9328 (
            .O(N__42347),
            .I(N__42341));
    InMux I__9327 (
            .O(N__42346),
            .I(N__42341));
    LocalMux I__9326 (
            .O(N__42341),
            .I(N__42337));
    InMux I__9325 (
            .O(N__42340),
            .I(N__42334));
    Span4Mux_h I__9324 (
            .O(N__42337),
            .I(N__42331));
    LocalMux I__9323 (
            .O(N__42334),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__9322 (
            .O(N__42331),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__9321 (
            .O(N__42326),
            .I(N__42323));
    LocalMux I__9320 (
            .O(N__42323),
            .I(N__42319));
    InMux I__9319 (
            .O(N__42322),
            .I(N__42314));
    Span4Mux_v I__9318 (
            .O(N__42319),
            .I(N__42311));
    InMux I__9317 (
            .O(N__42318),
            .I(N__42308));
    InMux I__9316 (
            .O(N__42317),
            .I(N__42305));
    LocalMux I__9315 (
            .O(N__42314),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__9314 (
            .O(N__42311),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    LocalMux I__9313 (
            .O(N__42308),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    LocalMux I__9312 (
            .O(N__42305),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__9311 (
            .O(N__42296),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__9310 (
            .O(N__42293),
            .I(N__42290));
    InMux I__9309 (
            .O(N__42290),
            .I(N__42286));
    InMux I__9308 (
            .O(N__42289),
            .I(N__42283));
    LocalMux I__9307 (
            .O(N__42286),
            .I(N__42277));
    LocalMux I__9306 (
            .O(N__42283),
            .I(N__42277));
    InMux I__9305 (
            .O(N__42282),
            .I(N__42274));
    Span4Mux_h I__9304 (
            .O(N__42277),
            .I(N__42271));
    LocalMux I__9303 (
            .O(N__42274),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__9302 (
            .O(N__42271),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__9301 (
            .O(N__42266),
            .I(N__42263));
    LocalMux I__9300 (
            .O(N__42263),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__9299 (
            .O(N__42260),
            .I(N__42257));
    LocalMux I__9298 (
            .O(N__42257),
            .I(N__42254));
    Odrv4 I__9297 (
            .O(N__42254),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__9296 (
            .O(N__42251),
            .I(N__42248));
    LocalMux I__9295 (
            .O(N__42248),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__9294 (
            .O(N__42245),
            .I(N__42242));
    LocalMux I__9293 (
            .O(N__42242),
            .I(N__42239));
    Odrv4 I__9292 (
            .O(N__42239),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__9291 (
            .O(N__42236),
            .I(N__42233));
    LocalMux I__9290 (
            .O(N__42233),
            .I(N__42230));
    Odrv4 I__9289 (
            .O(N__42230),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__9288 (
            .O(N__42227),
            .I(N__42224));
    LocalMux I__9287 (
            .O(N__42224),
            .I(N__42221));
    Span4Mux_v I__9286 (
            .O(N__42221),
            .I(N__42218));
    Odrv4 I__9285 (
            .O(N__42218),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__9284 (
            .O(N__42215),
            .I(N__42212));
    LocalMux I__9283 (
            .O(N__42212),
            .I(N__42209));
    Odrv4 I__9282 (
            .O(N__42209),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__9281 (
            .O(N__42206),
            .I(N__42203));
    LocalMux I__9280 (
            .O(N__42203),
            .I(N__42200));
    Odrv4 I__9279 (
            .O(N__42200),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    CascadeMux I__9278 (
            .O(N__42197),
            .I(N__42194));
    InMux I__9277 (
            .O(N__42194),
            .I(N__42191));
    LocalMux I__9276 (
            .O(N__42191),
            .I(N__42188));
    Odrv4 I__9275 (
            .O(N__42188),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    CascadeMux I__9274 (
            .O(N__42185),
            .I(N__42182));
    InMux I__9273 (
            .O(N__42182),
            .I(N__42179));
    LocalMux I__9272 (
            .O(N__42179),
            .I(N__42174));
    InMux I__9271 (
            .O(N__42178),
            .I(N__42171));
    InMux I__9270 (
            .O(N__42177),
            .I(N__42168));
    Odrv12 I__9269 (
            .O(N__42174),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__9268 (
            .O(N__42171),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__9267 (
            .O(N__42168),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__9266 (
            .O(N__42161),
            .I(N__42158));
    InMux I__9265 (
            .O(N__42158),
            .I(N__42155));
    LocalMux I__9264 (
            .O(N__42155),
            .I(N__42152));
    Odrv4 I__9263 (
            .O(N__42152),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    CascadeMux I__9262 (
            .O(N__42149),
            .I(N__42146));
    InMux I__9261 (
            .O(N__42146),
            .I(N__42143));
    LocalMux I__9260 (
            .O(N__42143),
            .I(N__42140));
    Odrv4 I__9259 (
            .O(N__42140),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__9258 (
            .O(N__42137),
            .I(N__42134));
    LocalMux I__9257 (
            .O(N__42134),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    CascadeMux I__9256 (
            .O(N__42131),
            .I(N__42128));
    InMux I__9255 (
            .O(N__42128),
            .I(N__42125));
    LocalMux I__9254 (
            .O(N__42125),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__9253 (
            .O(N__42122),
            .I(N__42119));
    LocalMux I__9252 (
            .O(N__42119),
            .I(N__42116));
    Odrv12 I__9251 (
            .O(N__42116),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__9250 (
            .O(N__42113),
            .I(N__42110));
    LocalMux I__9249 (
            .O(N__42110),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__9248 (
            .O(N__42107),
            .I(N__42104));
    LocalMux I__9247 (
            .O(N__42104),
            .I(N__42101));
    Odrv4 I__9246 (
            .O(N__42101),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__9245 (
            .O(N__42098),
            .I(N__42095));
    LocalMux I__9244 (
            .O(N__42095),
            .I(N__42092));
    Odrv4 I__9243 (
            .O(N__42092),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__9242 (
            .O(N__42089),
            .I(N__42086));
    LocalMux I__9241 (
            .O(N__42086),
            .I(N__42083));
    Odrv4 I__9240 (
            .O(N__42083),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__9239 (
            .O(N__42080),
            .I(N__42075));
    InMux I__9238 (
            .O(N__42079),
            .I(N__42072));
    InMux I__9237 (
            .O(N__42078),
            .I(N__42069));
    LocalMux I__9236 (
            .O(N__42075),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9235 (
            .O(N__42072),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9234 (
            .O(N__42069),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__9233 (
            .O(N__42062),
            .I(N__42059));
    LocalMux I__9232 (
            .O(N__42059),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    InMux I__9231 (
            .O(N__42056),
            .I(N__42053));
    LocalMux I__9230 (
            .O(N__42053),
            .I(N__42048));
    InMux I__9229 (
            .O(N__42052),
            .I(N__42045));
    InMux I__9228 (
            .O(N__42051),
            .I(N__42042));
    Odrv4 I__9227 (
            .O(N__42048),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__9226 (
            .O(N__42045),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__9225 (
            .O(N__42042),
            .I(\current_shift_inst.un4_control_input1_25 ));
    CascadeMux I__9224 (
            .O(N__42035),
            .I(N__42032));
    InMux I__9223 (
            .O(N__42032),
            .I(N__42029));
    LocalMux I__9222 (
            .O(N__42029),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__9221 (
            .O(N__42026),
            .I(N__42023));
    LocalMux I__9220 (
            .O(N__42023),
            .I(N__42018));
    CascadeMux I__9219 (
            .O(N__42022),
            .I(N__42015));
    InMux I__9218 (
            .O(N__42021),
            .I(N__42012));
    Span4Mux_v I__9217 (
            .O(N__42018),
            .I(N__42009));
    InMux I__9216 (
            .O(N__42015),
            .I(N__42006));
    LocalMux I__9215 (
            .O(N__42012),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__9214 (
            .O(N__42009),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__9213 (
            .O(N__42006),
            .I(\current_shift_inst.un4_control_input1_27 ));
    CascadeMux I__9212 (
            .O(N__41999),
            .I(N__41996));
    InMux I__9211 (
            .O(N__41996),
            .I(N__41993));
    LocalMux I__9210 (
            .O(N__41993),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__9209 (
            .O(N__41990),
            .I(N__41987));
    LocalMux I__9208 (
            .O(N__41987),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    CascadeMux I__9207 (
            .O(N__41984),
            .I(N__41979));
    InMux I__9206 (
            .O(N__41983),
            .I(N__41976));
    InMux I__9205 (
            .O(N__41982),
            .I(N__41973));
    InMux I__9204 (
            .O(N__41979),
            .I(N__41970));
    LocalMux I__9203 (
            .O(N__41976),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__9202 (
            .O(N__41973),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__9201 (
            .O(N__41970),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__9200 (
            .O(N__41963),
            .I(N__41960));
    LocalMux I__9199 (
            .O(N__41960),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    InMux I__9198 (
            .O(N__41957),
            .I(N__41954));
    LocalMux I__9197 (
            .O(N__41954),
            .I(N__41951));
    Odrv4 I__9196 (
            .O(N__41951),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__9195 (
            .O(N__41948),
            .I(N__41943));
    InMux I__9194 (
            .O(N__41947),
            .I(N__41940));
    InMux I__9193 (
            .O(N__41946),
            .I(N__41937));
    LocalMux I__9192 (
            .O(N__41943),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__9191 (
            .O(N__41940),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__9190 (
            .O(N__41937),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__9189 (
            .O(N__41930),
            .I(N__41927));
    LocalMux I__9188 (
            .O(N__41927),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__9187 (
            .O(N__41924),
            .I(N__41921));
    InMux I__9186 (
            .O(N__41921),
            .I(N__41918));
    LocalMux I__9185 (
            .O(N__41918),
            .I(N__41913));
    InMux I__9184 (
            .O(N__41917),
            .I(N__41910));
    InMux I__9183 (
            .O(N__41916),
            .I(N__41907));
    Odrv4 I__9182 (
            .O(N__41913),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__9181 (
            .O(N__41910),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__9180 (
            .O(N__41907),
            .I(\current_shift_inst.un4_control_input1_19 ));
    CascadeMux I__9179 (
            .O(N__41900),
            .I(N__41897));
    InMux I__9178 (
            .O(N__41897),
            .I(N__41894));
    LocalMux I__9177 (
            .O(N__41894),
            .I(N__41891));
    Odrv4 I__9176 (
            .O(N__41891),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__9175 (
            .O(N__41888),
            .I(N__41885));
    InMux I__9174 (
            .O(N__41885),
            .I(N__41882));
    LocalMux I__9173 (
            .O(N__41882),
            .I(N__41879));
    Odrv4 I__9172 (
            .O(N__41879),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__9171 (
            .O(N__41876),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__9170 (
            .O(N__41873),
            .I(N__41858));
    InMux I__9169 (
            .O(N__41872),
            .I(N__41855));
    InMux I__9168 (
            .O(N__41871),
            .I(N__41838));
    InMux I__9167 (
            .O(N__41870),
            .I(N__41838));
    InMux I__9166 (
            .O(N__41869),
            .I(N__41838));
    InMux I__9165 (
            .O(N__41868),
            .I(N__41838));
    InMux I__9164 (
            .O(N__41867),
            .I(N__41838));
    InMux I__9163 (
            .O(N__41866),
            .I(N__41838));
    InMux I__9162 (
            .O(N__41865),
            .I(N__41838));
    InMux I__9161 (
            .O(N__41864),
            .I(N__41838));
    CascadeMux I__9160 (
            .O(N__41863),
            .I(N__41834));
    InMux I__9159 (
            .O(N__41862),
            .I(N__41831));
    InMux I__9158 (
            .O(N__41861),
            .I(N__41828));
    LocalMux I__9157 (
            .O(N__41858),
            .I(N__41815));
    LocalMux I__9156 (
            .O(N__41855),
            .I(N__41815));
    LocalMux I__9155 (
            .O(N__41838),
            .I(N__41815));
    InMux I__9154 (
            .O(N__41837),
            .I(N__41812));
    InMux I__9153 (
            .O(N__41834),
            .I(N__41797));
    LocalMux I__9152 (
            .O(N__41831),
            .I(N__41792));
    LocalMux I__9151 (
            .O(N__41828),
            .I(N__41792));
    InMux I__9150 (
            .O(N__41827),
            .I(N__41789));
    InMux I__9149 (
            .O(N__41826),
            .I(N__41778));
    InMux I__9148 (
            .O(N__41825),
            .I(N__41778));
    InMux I__9147 (
            .O(N__41824),
            .I(N__41778));
    InMux I__9146 (
            .O(N__41823),
            .I(N__41778));
    InMux I__9145 (
            .O(N__41822),
            .I(N__41778));
    Span4Mux_v I__9144 (
            .O(N__41815),
            .I(N__41773));
    LocalMux I__9143 (
            .O(N__41812),
            .I(N__41773));
    InMux I__9142 (
            .O(N__41811),
            .I(N__41756));
    InMux I__9141 (
            .O(N__41810),
            .I(N__41756));
    InMux I__9140 (
            .O(N__41809),
            .I(N__41756));
    InMux I__9139 (
            .O(N__41808),
            .I(N__41756));
    InMux I__9138 (
            .O(N__41807),
            .I(N__41756));
    InMux I__9137 (
            .O(N__41806),
            .I(N__41756));
    InMux I__9136 (
            .O(N__41805),
            .I(N__41756));
    InMux I__9135 (
            .O(N__41804),
            .I(N__41756));
    InMux I__9134 (
            .O(N__41803),
            .I(N__41747));
    InMux I__9133 (
            .O(N__41802),
            .I(N__41747));
    InMux I__9132 (
            .O(N__41801),
            .I(N__41747));
    InMux I__9131 (
            .O(N__41800),
            .I(N__41747));
    LocalMux I__9130 (
            .O(N__41797),
            .I(N__41744));
    Span4Mux_v I__9129 (
            .O(N__41792),
            .I(N__41737));
    LocalMux I__9128 (
            .O(N__41789),
            .I(N__41737));
    LocalMux I__9127 (
            .O(N__41778),
            .I(N__41737));
    Span4Mux_h I__9126 (
            .O(N__41773),
            .I(N__41734));
    LocalMux I__9125 (
            .O(N__41756),
            .I(N__41729));
    LocalMux I__9124 (
            .O(N__41747),
            .I(N__41729));
    Odrv4 I__9123 (
            .O(N__41744),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__9122 (
            .O(N__41737),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__9121 (
            .O(N__41734),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv12 I__9120 (
            .O(N__41729),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__9119 (
            .O(N__41720),
            .I(N__41717));
    LocalMux I__9118 (
            .O(N__41717),
            .I(N__41712));
    InMux I__9117 (
            .O(N__41716),
            .I(N__41709));
    InMux I__9116 (
            .O(N__41715),
            .I(N__41706));
    Odrv4 I__9115 (
            .O(N__41712),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__9114 (
            .O(N__41709),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__9113 (
            .O(N__41706),
            .I(\current_shift_inst.un4_control_input1_29 ));
    CascadeMux I__9112 (
            .O(N__41699),
            .I(N__41696));
    InMux I__9111 (
            .O(N__41696),
            .I(N__41693));
    LocalMux I__9110 (
            .O(N__41693),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__9109 (
            .O(N__41690),
            .I(N__41687));
    LocalMux I__9108 (
            .O(N__41687),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__9107 (
            .O(N__41684),
            .I(N__41681));
    LocalMux I__9106 (
            .O(N__41681),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__9105 (
            .O(N__41678),
            .I(N__41675));
    InMux I__9104 (
            .O(N__41675),
            .I(N__41672));
    LocalMux I__9103 (
            .O(N__41672),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__9102 (
            .O(N__41669),
            .I(N__41666));
    InMux I__9101 (
            .O(N__41666),
            .I(N__41663));
    LocalMux I__9100 (
            .O(N__41663),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    CascadeMux I__9099 (
            .O(N__41660),
            .I(N__41657));
    InMux I__9098 (
            .O(N__41657),
            .I(N__41654));
    LocalMux I__9097 (
            .O(N__41654),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__9096 (
            .O(N__41651),
            .I(N__41648));
    InMux I__9095 (
            .O(N__41648),
            .I(N__41645));
    LocalMux I__9094 (
            .O(N__41645),
            .I(N__41642));
    Span4Mux_h I__9093 (
            .O(N__41642),
            .I(N__41639));
    Odrv4 I__9092 (
            .O(N__41639),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    CascadeMux I__9091 (
            .O(N__41636),
            .I(N__41633));
    InMux I__9090 (
            .O(N__41633),
            .I(N__41630));
    LocalMux I__9089 (
            .O(N__41630),
            .I(N__41627));
    Odrv4 I__9088 (
            .O(N__41627),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    InMux I__9087 (
            .O(N__41624),
            .I(N__41621));
    LocalMux I__9086 (
            .O(N__41621),
            .I(N__41618));
    Span4Mux_h I__9085 (
            .O(N__41618),
            .I(N__41615));
    Odrv4 I__9084 (
            .O(N__41615),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    CascadeMux I__9083 (
            .O(N__41612),
            .I(N__41609));
    InMux I__9082 (
            .O(N__41609),
            .I(N__41606));
    LocalMux I__9081 (
            .O(N__41606),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__9080 (
            .O(N__41603),
            .I(N__41600));
    LocalMux I__9079 (
            .O(N__41600),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__9078 (
            .O(N__41597),
            .I(N__41594));
    InMux I__9077 (
            .O(N__41594),
            .I(N__41591));
    LocalMux I__9076 (
            .O(N__41591),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__9075 (
            .O(N__41588),
            .I(N__41585));
    LocalMux I__9074 (
            .O(N__41585),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__9073 (
            .O(N__41582),
            .I(N__41579));
    InMux I__9072 (
            .O(N__41579),
            .I(N__41576));
    LocalMux I__9071 (
            .O(N__41576),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__9070 (
            .O(N__41573),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__9069 (
            .O(N__41570),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__9068 (
            .O(N__41567),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__9067 (
            .O(N__41564),
            .I(N__41526));
    InMux I__9066 (
            .O(N__41563),
            .I(N__41526));
    InMux I__9065 (
            .O(N__41562),
            .I(N__41526));
    InMux I__9064 (
            .O(N__41561),
            .I(N__41526));
    InMux I__9063 (
            .O(N__41560),
            .I(N__41517));
    InMux I__9062 (
            .O(N__41559),
            .I(N__41517));
    InMux I__9061 (
            .O(N__41558),
            .I(N__41517));
    InMux I__9060 (
            .O(N__41557),
            .I(N__41517));
    InMux I__9059 (
            .O(N__41556),
            .I(N__41508));
    InMux I__9058 (
            .O(N__41555),
            .I(N__41508));
    InMux I__9057 (
            .O(N__41554),
            .I(N__41508));
    InMux I__9056 (
            .O(N__41553),
            .I(N__41508));
    InMux I__9055 (
            .O(N__41552),
            .I(N__41499));
    InMux I__9054 (
            .O(N__41551),
            .I(N__41499));
    InMux I__9053 (
            .O(N__41550),
            .I(N__41499));
    InMux I__9052 (
            .O(N__41549),
            .I(N__41499));
    InMux I__9051 (
            .O(N__41548),
            .I(N__41490));
    InMux I__9050 (
            .O(N__41547),
            .I(N__41490));
    InMux I__9049 (
            .O(N__41546),
            .I(N__41490));
    InMux I__9048 (
            .O(N__41545),
            .I(N__41490));
    InMux I__9047 (
            .O(N__41544),
            .I(N__41481));
    InMux I__9046 (
            .O(N__41543),
            .I(N__41481));
    InMux I__9045 (
            .O(N__41542),
            .I(N__41481));
    InMux I__9044 (
            .O(N__41541),
            .I(N__41481));
    InMux I__9043 (
            .O(N__41540),
            .I(N__41476));
    InMux I__9042 (
            .O(N__41539),
            .I(N__41476));
    InMux I__9041 (
            .O(N__41538),
            .I(N__41467));
    InMux I__9040 (
            .O(N__41537),
            .I(N__41467));
    InMux I__9039 (
            .O(N__41536),
            .I(N__41467));
    InMux I__9038 (
            .O(N__41535),
            .I(N__41467));
    LocalMux I__9037 (
            .O(N__41526),
            .I(N__41462));
    LocalMux I__9036 (
            .O(N__41517),
            .I(N__41462));
    LocalMux I__9035 (
            .O(N__41508),
            .I(N__41459));
    LocalMux I__9034 (
            .O(N__41499),
            .I(N__41448));
    LocalMux I__9033 (
            .O(N__41490),
            .I(N__41448));
    LocalMux I__9032 (
            .O(N__41481),
            .I(N__41448));
    LocalMux I__9031 (
            .O(N__41476),
            .I(N__41448));
    LocalMux I__9030 (
            .O(N__41467),
            .I(N__41448));
    Span4Mux_v I__9029 (
            .O(N__41462),
            .I(N__41441));
    Span4Mux_h I__9028 (
            .O(N__41459),
            .I(N__41441));
    Span4Mux_v I__9027 (
            .O(N__41448),
            .I(N__41441));
    Span4Mux_h I__9026 (
            .O(N__41441),
            .I(N__41438));
    Odrv4 I__9025 (
            .O(N__41438),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__9024 (
            .O(N__41435),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CEMux I__9023 (
            .O(N__41432),
            .I(N__41427));
    CEMux I__9022 (
            .O(N__41431),
            .I(N__41424));
    CEMux I__9021 (
            .O(N__41430),
            .I(N__41421));
    LocalMux I__9020 (
            .O(N__41427),
            .I(N__41417));
    LocalMux I__9019 (
            .O(N__41424),
            .I(N__41414));
    LocalMux I__9018 (
            .O(N__41421),
            .I(N__41411));
    CEMux I__9017 (
            .O(N__41420),
            .I(N__41408));
    Span4Mux_h I__9016 (
            .O(N__41417),
            .I(N__41405));
    Span4Mux_h I__9015 (
            .O(N__41414),
            .I(N__41402));
    Span4Mux_v I__9014 (
            .O(N__41411),
            .I(N__41399));
    LocalMux I__9013 (
            .O(N__41408),
            .I(N__41396));
    Span4Mux_v I__9012 (
            .O(N__41405),
            .I(N__41393));
    Span4Mux_h I__9011 (
            .O(N__41402),
            .I(N__41390));
    Span4Mux_h I__9010 (
            .O(N__41399),
            .I(N__41385));
    Span4Mux_v I__9009 (
            .O(N__41396),
            .I(N__41385));
    Odrv4 I__9008 (
            .O(N__41393),
            .I(\delay_measurement_inst.delay_hc_timer.N_164_i ));
    Odrv4 I__9007 (
            .O(N__41390),
            .I(\delay_measurement_inst.delay_hc_timer.N_164_i ));
    Odrv4 I__9006 (
            .O(N__41385),
            .I(\delay_measurement_inst.delay_hc_timer.N_164_i ));
    CascadeMux I__9005 (
            .O(N__41378),
            .I(N__41375));
    InMux I__9004 (
            .O(N__41375),
            .I(N__41372));
    LocalMux I__9003 (
            .O(N__41372),
            .I(N__41369));
    Span4Mux_v I__9002 (
            .O(N__41369),
            .I(N__41366));
    Odrv4 I__9001 (
            .O(N__41366),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__9000 (
            .O(N__41363),
            .I(N__41360));
    LocalMux I__8999 (
            .O(N__41360),
            .I(N__41357));
    Span4Mux_h I__8998 (
            .O(N__41357),
            .I(N__41354));
    Odrv4 I__8997 (
            .O(N__41354),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    CascadeMux I__8996 (
            .O(N__41351),
            .I(N__41348));
    InMux I__8995 (
            .O(N__41348),
            .I(N__41345));
    LocalMux I__8994 (
            .O(N__41345),
            .I(N__41342));
    Odrv12 I__8993 (
            .O(N__41342),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    InMux I__8992 (
            .O(N__41339),
            .I(N__41335));
    InMux I__8991 (
            .O(N__41338),
            .I(N__41332));
    LocalMux I__8990 (
            .O(N__41335),
            .I(N__41328));
    LocalMux I__8989 (
            .O(N__41332),
            .I(N__41325));
    InMux I__8988 (
            .O(N__41331),
            .I(N__41322));
    Odrv4 I__8987 (
            .O(N__41328),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv12 I__8986 (
            .O(N__41325),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__8985 (
            .O(N__41322),
            .I(\current_shift_inst.un4_control_input1_5 ));
    CascadeMux I__8984 (
            .O(N__41315),
            .I(N__41312));
    InMux I__8983 (
            .O(N__41312),
            .I(N__41309));
    LocalMux I__8982 (
            .O(N__41309),
            .I(N__41306));
    Span4Mux_h I__8981 (
            .O(N__41306),
            .I(N__41303));
    Odrv4 I__8980 (
            .O(N__41303),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ));
    CascadeMux I__8979 (
            .O(N__41300),
            .I(N__41297));
    InMux I__8978 (
            .O(N__41297),
            .I(N__41294));
    LocalMux I__8977 (
            .O(N__41294),
            .I(N__41291));
    Span4Mux_h I__8976 (
            .O(N__41291),
            .I(N__41288));
    Odrv4 I__8975 (
            .O(N__41288),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    InMux I__8974 (
            .O(N__41285),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__8973 (
            .O(N__41282),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__8972 (
            .O(N__41279),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__8971 (
            .O(N__41276),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__8970 (
            .O(N__41273),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__8969 (
            .O(N__41270),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__8968 (
            .O(N__41267),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__8967 (
            .O(N__41264),
            .I(bfn_17_13_0_));
    InMux I__8966 (
            .O(N__41261),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__8965 (
            .O(N__41258),
            .I(bfn_17_11_0_));
    InMux I__8964 (
            .O(N__41255),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__8963 (
            .O(N__41252),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__8962 (
            .O(N__41249),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__8961 (
            .O(N__41246),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__8960 (
            .O(N__41243),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__8959 (
            .O(N__41240),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__8958 (
            .O(N__41237),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__8957 (
            .O(N__41234),
            .I(bfn_17_12_0_));
    CascadeMux I__8956 (
            .O(N__41231),
            .I(elapsed_time_ns_1_RNI02CN9_0_13_cascade_));
    InMux I__8955 (
            .O(N__41228),
            .I(N__41225));
    LocalMux I__8954 (
            .O(N__41225),
            .I(N__41222));
    Span4Mux_h I__8953 (
            .O(N__41222),
            .I(N__41219));
    Odrv4 I__8952 (
            .O(N__41219),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__8951 (
            .O(N__41216),
            .I(bfn_17_10_0_));
    InMux I__8950 (
            .O(N__41213),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__8949 (
            .O(N__41210),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__8948 (
            .O(N__41207),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__8947 (
            .O(N__41204),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__8946 (
            .O(N__41201),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__8945 (
            .O(N__41198),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__8944 (
            .O(N__41195),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__8943 (
            .O(N__41192),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ));
    InMux I__8942 (
            .O(N__41189),
            .I(N__41186));
    LocalMux I__8941 (
            .O(N__41186),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    InMux I__8940 (
            .O(N__41183),
            .I(N__41180));
    LocalMux I__8939 (
            .O(N__41180),
            .I(N__41177));
    Odrv4 I__8938 (
            .O(N__41177),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    InMux I__8937 (
            .O(N__41174),
            .I(N__41171));
    LocalMux I__8936 (
            .O(N__41171),
            .I(N__41167));
    InMux I__8935 (
            .O(N__41170),
            .I(N__41163));
    Span4Mux_v I__8934 (
            .O(N__41167),
            .I(N__41160));
    InMux I__8933 (
            .O(N__41166),
            .I(N__41157));
    LocalMux I__8932 (
            .O(N__41163),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__8931 (
            .O(N__41160),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    LocalMux I__8930 (
            .O(N__41157),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    CascadeMux I__8929 (
            .O(N__41150),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_ ));
    InMux I__8928 (
            .O(N__41147),
            .I(N__41144));
    LocalMux I__8927 (
            .O(N__41144),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    CascadeMux I__8926 (
            .O(N__41141),
            .I(N__41138));
    InMux I__8925 (
            .O(N__41138),
            .I(N__41135));
    LocalMux I__8924 (
            .O(N__41135),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    InMux I__8923 (
            .O(N__41132),
            .I(N__41129));
    LocalMux I__8922 (
            .O(N__41129),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ));
    InMux I__8921 (
            .O(N__41126),
            .I(N__41123));
    LocalMux I__8920 (
            .O(N__41123),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    InMux I__8919 (
            .O(N__41120),
            .I(N__41116));
    InMux I__8918 (
            .O(N__41119),
            .I(N__41113));
    LocalMux I__8917 (
            .O(N__41116),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__8916 (
            .O(N__41113),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    InMux I__8915 (
            .O(N__41108),
            .I(N__41105));
    LocalMux I__8914 (
            .O(N__41105),
            .I(N__41102));
    Span4Mux_h I__8913 (
            .O(N__41102),
            .I(N__41099));
    Odrv4 I__8912 (
            .O(N__41099),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__8911 (
            .O(N__41096),
            .I(N__41093));
    LocalMux I__8910 (
            .O(N__41093),
            .I(N__41090));
    Span4Mux_v I__8909 (
            .O(N__41090),
            .I(N__41086));
    InMux I__8908 (
            .O(N__41089),
            .I(N__41083));
    Odrv4 I__8907 (
            .O(N__41086),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    LocalMux I__8906 (
            .O(N__41083),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    CascadeMux I__8905 (
            .O(N__41078),
            .I(elapsed_time_ns_1_RNITUBN9_0_10_cascade_));
    InMux I__8904 (
            .O(N__41075),
            .I(N__41072));
    LocalMux I__8903 (
            .O(N__41072),
            .I(N__41069));
    Span4Mux_v I__8902 (
            .O(N__41069),
            .I(N__41066));
    Odrv4 I__8901 (
            .O(N__41066),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__8900 (
            .O(N__41063),
            .I(N__41060));
    LocalMux I__8899 (
            .O(N__41060),
            .I(N__41056));
    InMux I__8898 (
            .O(N__41059),
            .I(N__41052));
    Span4Mux_v I__8897 (
            .O(N__41056),
            .I(N__41049));
    InMux I__8896 (
            .O(N__41055),
            .I(N__41046));
    LocalMux I__8895 (
            .O(N__41052),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv4 I__8894 (
            .O(N__41049),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    LocalMux I__8893 (
            .O(N__41046),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    InMux I__8892 (
            .O(N__41039),
            .I(N__41036));
    LocalMux I__8891 (
            .O(N__41036),
            .I(N__41033));
    Span4Mux_h I__8890 (
            .O(N__41033),
            .I(N__41030));
    Odrv4 I__8889 (
            .O(N__41030),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__8888 (
            .O(N__41027),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ));
    InMux I__8887 (
            .O(N__41024),
            .I(N__41021));
    LocalMux I__8886 (
            .O(N__41021),
            .I(N__41018));
    Span4Mux_h I__8885 (
            .O(N__41018),
            .I(N__41015));
    Odrv4 I__8884 (
            .O(N__41015),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    CascadeMux I__8883 (
            .O(N__41012),
            .I(N__41009));
    InMux I__8882 (
            .O(N__41009),
            .I(N__41005));
    InMux I__8881 (
            .O(N__41008),
            .I(N__41002));
    LocalMux I__8880 (
            .O(N__41005),
            .I(N__40998));
    LocalMux I__8879 (
            .O(N__41002),
            .I(N__40995));
    InMux I__8878 (
            .O(N__41001),
            .I(N__40992));
    Odrv4 I__8877 (
            .O(N__40998),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv12 I__8876 (
            .O(N__40995),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    LocalMux I__8875 (
            .O(N__40992),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__8874 (
            .O(N__40985),
            .I(N__40982));
    InMux I__8873 (
            .O(N__40982),
            .I(N__40979));
    LocalMux I__8872 (
            .O(N__40979),
            .I(N__40976));
    Odrv12 I__8871 (
            .O(N__40976),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    InMux I__8870 (
            .O(N__40973),
            .I(N__40969));
    InMux I__8869 (
            .O(N__40972),
            .I(N__40966));
    LocalMux I__8868 (
            .O(N__40969),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    LocalMux I__8867 (
            .O(N__40966),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__8866 (
            .O(N__40961),
            .I(N__40957));
    InMux I__8865 (
            .O(N__40960),
            .I(N__40954));
    LocalMux I__8864 (
            .O(N__40957),
            .I(N__40948));
    LocalMux I__8863 (
            .O(N__40954),
            .I(N__40948));
    InMux I__8862 (
            .O(N__40953),
            .I(N__40945));
    Span4Mux_h I__8861 (
            .O(N__40948),
            .I(N__40942));
    LocalMux I__8860 (
            .O(N__40945),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__8859 (
            .O(N__40942),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__8858 (
            .O(N__40937),
            .I(N__40933));
    InMux I__8857 (
            .O(N__40936),
            .I(N__40928));
    InMux I__8856 (
            .O(N__40933),
            .I(N__40928));
    LocalMux I__8855 (
            .O(N__40928),
            .I(N__40924));
    InMux I__8854 (
            .O(N__40927),
            .I(N__40921));
    Span4Mux_h I__8853 (
            .O(N__40924),
            .I(N__40918));
    LocalMux I__8852 (
            .O(N__40921),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__8851 (
            .O(N__40918),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__8850 (
            .O(N__40913),
            .I(N__40910));
    LocalMux I__8849 (
            .O(N__40910),
            .I(N__40907));
    Span4Mux_h I__8848 (
            .O(N__40907),
            .I(N__40904));
    Odrv4 I__8847 (
            .O(N__40904),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__8846 (
            .O(N__40901),
            .I(N__40898));
    LocalMux I__8845 (
            .O(N__40898),
            .I(N__40895));
    Span4Mux_v I__8844 (
            .O(N__40895),
            .I(N__40891));
    InMux I__8843 (
            .O(N__40894),
            .I(N__40888));
    Odrv4 I__8842 (
            .O(N__40891),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    LocalMux I__8841 (
            .O(N__40888),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    CascadeMux I__8840 (
            .O(N__40883),
            .I(elapsed_time_ns_1_RNI46CN9_0_17_cascade_));
    CascadeMux I__8839 (
            .O(N__40880),
            .I(N__40877));
    InMux I__8838 (
            .O(N__40877),
            .I(N__40871));
    InMux I__8837 (
            .O(N__40876),
            .I(N__40871));
    LocalMux I__8836 (
            .O(N__40871),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__8835 (
            .O(N__40868),
            .I(N__40865));
    LocalMux I__8834 (
            .O(N__40865),
            .I(N__40861));
    InMux I__8833 (
            .O(N__40864),
            .I(N__40857));
    Span4Mux_v I__8832 (
            .O(N__40861),
            .I(N__40854));
    InMux I__8831 (
            .O(N__40860),
            .I(N__40851));
    LocalMux I__8830 (
            .O(N__40857),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__8829 (
            .O(N__40854),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    LocalMux I__8828 (
            .O(N__40851),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__8827 (
            .O(N__40844),
            .I(N__40840));
    InMux I__8826 (
            .O(N__40843),
            .I(N__40837));
    LocalMux I__8825 (
            .O(N__40840),
            .I(N__40831));
    LocalMux I__8824 (
            .O(N__40837),
            .I(N__40831));
    InMux I__8823 (
            .O(N__40836),
            .I(N__40828));
    Span4Mux_v I__8822 (
            .O(N__40831),
            .I(N__40825));
    LocalMux I__8821 (
            .O(N__40828),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    Odrv4 I__8820 (
            .O(N__40825),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    InMux I__8819 (
            .O(N__40820),
            .I(N__40817));
    LocalMux I__8818 (
            .O(N__40817),
            .I(N__40814));
    Span4Mux_v I__8817 (
            .O(N__40814),
            .I(N__40811));
    Odrv4 I__8816 (
            .O(N__40811),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__8815 (
            .O(N__40808),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__8814 (
            .O(N__40805),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__8813 (
            .O(N__40802),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__8812 (
            .O(N__40799),
            .I(bfn_16_20_0_));
    InMux I__8811 (
            .O(N__40796),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__8810 (
            .O(N__40793),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__8809 (
            .O(N__40790),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__8808 (
            .O(N__40787),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__8807 (
            .O(N__40784),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__8806 (
            .O(N__40781),
            .I(N__40778));
    LocalMux I__8805 (
            .O(N__40778),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__8804 (
            .O(N__40775),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__8803 (
            .O(N__40772),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__8802 (
            .O(N__40769),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__8801 (
            .O(N__40766),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__8800 (
            .O(N__40763),
            .I(bfn_16_19_0_));
    InMux I__8799 (
            .O(N__40760),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__8798 (
            .O(N__40757),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__8797 (
            .O(N__40754),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__8796 (
            .O(N__40751),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__8795 (
            .O(N__40748),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__8794 (
            .O(N__40745),
            .I(N__40742));
    LocalMux I__8793 (
            .O(N__40742),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__8792 (
            .O(N__40739),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    CascadeMux I__8791 (
            .O(N__40736),
            .I(N__40733));
    InMux I__8790 (
            .O(N__40733),
            .I(N__40729));
    InMux I__8789 (
            .O(N__40732),
            .I(N__40725));
    LocalMux I__8788 (
            .O(N__40729),
            .I(N__40722));
    InMux I__8787 (
            .O(N__40728),
            .I(N__40719));
    LocalMux I__8786 (
            .O(N__40725),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv12 I__8785 (
            .O(N__40722),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__8784 (
            .O(N__40719),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__8783 (
            .O(N__40712),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    CascadeMux I__8782 (
            .O(N__40709),
            .I(N__40705));
    InMux I__8781 (
            .O(N__40708),
            .I(N__40702));
    InMux I__8780 (
            .O(N__40705),
            .I(N__40699));
    LocalMux I__8779 (
            .O(N__40702),
            .I(N__40696));
    LocalMux I__8778 (
            .O(N__40699),
            .I(N__40692));
    Span4Mux_h I__8777 (
            .O(N__40696),
            .I(N__40689));
    InMux I__8776 (
            .O(N__40695),
            .I(N__40686));
    Odrv12 I__8775 (
            .O(N__40692),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__8774 (
            .O(N__40689),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__8773 (
            .O(N__40686),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__8772 (
            .O(N__40679),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__8771 (
            .O(N__40676),
            .I(N__40673));
    LocalMux I__8770 (
            .O(N__40673),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__8769 (
            .O(N__40670),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    CascadeMux I__8768 (
            .O(N__40667),
            .I(N__40663));
    InMux I__8767 (
            .O(N__40666),
            .I(N__40655));
    InMux I__8766 (
            .O(N__40663),
            .I(N__40655));
    InMux I__8765 (
            .O(N__40662),
            .I(N__40655));
    LocalMux I__8764 (
            .O(N__40655),
            .I(N__40652));
    Odrv4 I__8763 (
            .O(N__40652),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__8762 (
            .O(N__40649),
            .I(bfn_16_18_0_));
    InMux I__8761 (
            .O(N__40646),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__8760 (
            .O(N__40643),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__8759 (
            .O(N__40640),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__8758 (
            .O(N__40637),
            .I(N__40634));
    LocalMux I__8757 (
            .O(N__40634),
            .I(N__40631));
    Odrv4 I__8756 (
            .O(N__40631),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    InMux I__8755 (
            .O(N__40628),
            .I(N__40619));
    InMux I__8754 (
            .O(N__40627),
            .I(N__40619));
    InMux I__8753 (
            .O(N__40626),
            .I(N__40619));
    LocalMux I__8752 (
            .O(N__40619),
            .I(N__40616));
    Odrv4 I__8751 (
            .O(N__40616),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__8750 (
            .O(N__40613),
            .I(N__40610));
    LocalMux I__8749 (
            .O(N__40610),
            .I(N__40606));
    InMux I__8748 (
            .O(N__40609),
            .I(N__40603));
    Span4Mux_h I__8747 (
            .O(N__40606),
            .I(N__40599));
    LocalMux I__8746 (
            .O(N__40603),
            .I(N__40596));
    InMux I__8745 (
            .O(N__40602),
            .I(N__40593));
    Odrv4 I__8744 (
            .O(N__40599),
            .I(\current_shift_inst.un4_control_input1_3 ));
    Odrv12 I__8743 (
            .O(N__40596),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__8742 (
            .O(N__40593),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__8741 (
            .O(N__40586),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__8740 (
            .O(N__40583),
            .I(N__40577));
    InMux I__8739 (
            .O(N__40582),
            .I(N__40577));
    LocalMux I__8738 (
            .O(N__40577),
            .I(N__40574));
    Span4Mux_h I__8737 (
            .O(N__40574),
            .I(N__40570));
    InMux I__8736 (
            .O(N__40573),
            .I(N__40567));
    Odrv4 I__8735 (
            .O(N__40570),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__8734 (
            .O(N__40567),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__8733 (
            .O(N__40562),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__8732 (
            .O(N__40559),
            .I(N__40556));
    LocalMux I__8731 (
            .O(N__40556),
            .I(N__40553));
    Span4Mux_h I__8730 (
            .O(N__40553),
            .I(N__40550));
    Odrv4 I__8729 (
            .O(N__40550),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    InMux I__8728 (
            .O(N__40547),
            .I(N__40544));
    LocalMux I__8727 (
            .O(N__40544),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__8726 (
            .O(N__40541),
            .I(N__40538));
    LocalMux I__8725 (
            .O(N__40538),
            .I(N__40535));
    Span4Mux_h I__8724 (
            .O(N__40535),
            .I(N__40532));
    Odrv4 I__8723 (
            .O(N__40532),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    CascadeMux I__8722 (
            .O(N__40529),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    InMux I__8721 (
            .O(N__40526),
            .I(N__40523));
    LocalMux I__8720 (
            .O(N__40523),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ));
    InMux I__8719 (
            .O(N__40520),
            .I(N__40517));
    LocalMux I__8718 (
            .O(N__40517),
            .I(N__40514));
    Odrv4 I__8717 (
            .O(N__40514),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__8716 (
            .O(N__40511),
            .I(N__40508));
    LocalMux I__8715 (
            .O(N__40508),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    CascadeMux I__8714 (
            .O(N__40505),
            .I(N__40502));
    InMux I__8713 (
            .O(N__40502),
            .I(N__40499));
    LocalMux I__8712 (
            .O(N__40499),
            .I(N__40496));
    Span4Mux_h I__8711 (
            .O(N__40496),
            .I(N__40493));
    Odrv4 I__8710 (
            .O(N__40493),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__8709 (
            .O(N__40490),
            .I(N__40483));
    InMux I__8708 (
            .O(N__40489),
            .I(N__40483));
    CascadeMux I__8707 (
            .O(N__40488),
            .I(N__40480));
    LocalMux I__8706 (
            .O(N__40483),
            .I(N__40477));
    InMux I__8705 (
            .O(N__40480),
            .I(N__40474));
    Span4Mux_v I__8704 (
            .O(N__40477),
            .I(N__40470));
    LocalMux I__8703 (
            .O(N__40474),
            .I(N__40467));
    InMux I__8702 (
            .O(N__40473),
            .I(N__40464));
    Odrv4 I__8701 (
            .O(N__40470),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__8700 (
            .O(N__40467),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__8699 (
            .O(N__40464),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    InMux I__8698 (
            .O(N__40457),
            .I(N__40454));
    LocalMux I__8697 (
            .O(N__40454),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__8696 (
            .O(N__40451),
            .I(N__40447));
    InMux I__8695 (
            .O(N__40450),
            .I(N__40440));
    InMux I__8694 (
            .O(N__40447),
            .I(N__40440));
    InMux I__8693 (
            .O(N__40446),
            .I(N__40435));
    InMux I__8692 (
            .O(N__40445),
            .I(N__40435));
    LocalMux I__8691 (
            .O(N__40440),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__8690 (
            .O(N__40435),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__8689 (
            .O(N__40430),
            .I(N__40427));
    LocalMux I__8688 (
            .O(N__40427),
            .I(N__40424));
    Odrv4 I__8687 (
            .O(N__40424),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    InMux I__8686 (
            .O(N__40421),
            .I(N__40418));
    LocalMux I__8685 (
            .O(N__40418),
            .I(N__40414));
    InMux I__8684 (
            .O(N__40417),
            .I(N__40411));
    Odrv12 I__8683 (
            .O(N__40414),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    LocalMux I__8682 (
            .O(N__40411),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    InMux I__8681 (
            .O(N__40406),
            .I(N__40400));
    InMux I__8680 (
            .O(N__40405),
            .I(N__40400));
    LocalMux I__8679 (
            .O(N__40400),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    InMux I__8678 (
            .O(N__40397),
            .I(N__40394));
    LocalMux I__8677 (
            .O(N__40394),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    InMux I__8676 (
            .O(N__40391),
            .I(N__40388));
    LocalMux I__8675 (
            .O(N__40388),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    InMux I__8674 (
            .O(N__40385),
            .I(N__40382));
    LocalMux I__8673 (
            .O(N__40382),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__8672 (
            .O(N__40379),
            .I(N__40376));
    LocalMux I__8671 (
            .O(N__40376),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    CascadeMux I__8670 (
            .O(N__40373),
            .I(N__40370));
    InMux I__8669 (
            .O(N__40370),
            .I(N__40367));
    LocalMux I__8668 (
            .O(N__40367),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ));
    InMux I__8667 (
            .O(N__40364),
            .I(N__40361));
    LocalMux I__8666 (
            .O(N__40361),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    InMux I__8665 (
            .O(N__40358),
            .I(N__40355));
    LocalMux I__8664 (
            .O(N__40355),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    CascadeMux I__8663 (
            .O(N__40352),
            .I(N__40349));
    InMux I__8662 (
            .O(N__40349),
            .I(N__40346));
    LocalMux I__8661 (
            .O(N__40346),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    CascadeMux I__8660 (
            .O(N__40343),
            .I(N__40340));
    InMux I__8659 (
            .O(N__40340),
            .I(N__40337));
    LocalMux I__8658 (
            .O(N__40337),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    InMux I__8657 (
            .O(N__40334),
            .I(N__40328));
    InMux I__8656 (
            .O(N__40333),
            .I(N__40328));
    LocalMux I__8655 (
            .O(N__40328),
            .I(N__40324));
    InMux I__8654 (
            .O(N__40327),
            .I(N__40321));
    Span4Mux_h I__8653 (
            .O(N__40324),
            .I(N__40318));
    LocalMux I__8652 (
            .O(N__40321),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__8651 (
            .O(N__40318),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    CascadeMux I__8650 (
            .O(N__40313),
            .I(N__40310));
    InMux I__8649 (
            .O(N__40310),
            .I(N__40304));
    InMux I__8648 (
            .O(N__40309),
            .I(N__40304));
    LocalMux I__8647 (
            .O(N__40304),
            .I(N__40300));
    InMux I__8646 (
            .O(N__40303),
            .I(N__40297));
    Span4Mux_h I__8645 (
            .O(N__40300),
            .I(N__40294));
    LocalMux I__8644 (
            .O(N__40297),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__8643 (
            .O(N__40294),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__8642 (
            .O(N__40289),
            .I(N__40286));
    LocalMux I__8641 (
            .O(N__40286),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    InMux I__8640 (
            .O(N__40283),
            .I(N__40280));
    LocalMux I__8639 (
            .O(N__40280),
            .I(N__40277));
    Span4Mux_v I__8638 (
            .O(N__40277),
            .I(N__40273));
    InMux I__8637 (
            .O(N__40276),
            .I(N__40270));
    Odrv4 I__8636 (
            .O(N__40273),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__8635 (
            .O(N__40270),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    InMux I__8634 (
            .O(N__40265),
            .I(N__40259));
    InMux I__8633 (
            .O(N__40264),
            .I(N__40259));
    LocalMux I__8632 (
            .O(N__40259),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    InMux I__8631 (
            .O(N__40256),
            .I(N__40253));
    LocalMux I__8630 (
            .O(N__40253),
            .I(N__40250));
    Span4Mux_v I__8629 (
            .O(N__40250),
            .I(N__40245));
    InMux I__8628 (
            .O(N__40249),
            .I(N__40242));
    InMux I__8627 (
            .O(N__40248),
            .I(N__40239));
    Span4Mux_h I__8626 (
            .O(N__40245),
            .I(N__40234));
    LocalMux I__8625 (
            .O(N__40242),
            .I(N__40234));
    LocalMux I__8624 (
            .O(N__40239),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv4 I__8623 (
            .O(N__40234),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    CascadeMux I__8622 (
            .O(N__40229),
            .I(N__40226));
    InMux I__8621 (
            .O(N__40226),
            .I(N__40220));
    InMux I__8620 (
            .O(N__40225),
            .I(N__40220));
    LocalMux I__8619 (
            .O(N__40220),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    InMux I__8618 (
            .O(N__40217),
            .I(N__40212));
    InMux I__8617 (
            .O(N__40216),
            .I(N__40209));
    InMux I__8616 (
            .O(N__40215),
            .I(N__40206));
    LocalMux I__8615 (
            .O(N__40212),
            .I(N__40203));
    LocalMux I__8614 (
            .O(N__40209),
            .I(N__40200));
    LocalMux I__8613 (
            .O(N__40206),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    Odrv12 I__8612 (
            .O(N__40203),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    Odrv4 I__8611 (
            .O(N__40200),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    CascadeMux I__8610 (
            .O(N__40193),
            .I(N__40190));
    InMux I__8609 (
            .O(N__40190),
            .I(N__40187));
    LocalMux I__8608 (
            .O(N__40187),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__8607 (
            .O(N__40184),
            .I(N__40181));
    LocalMux I__8606 (
            .O(N__40181),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__8605 (
            .O(N__40178),
            .I(N__40175));
    InMux I__8604 (
            .O(N__40175),
            .I(N__40172));
    LocalMux I__8603 (
            .O(N__40172),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    CascadeMux I__8602 (
            .O(N__40169),
            .I(N__40165));
    InMux I__8601 (
            .O(N__40168),
            .I(N__40159));
    InMux I__8600 (
            .O(N__40165),
            .I(N__40159));
    InMux I__8599 (
            .O(N__40164),
            .I(N__40156));
    LocalMux I__8598 (
            .O(N__40159),
            .I(N__40153));
    LocalMux I__8597 (
            .O(N__40156),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__8596 (
            .O(N__40153),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    CascadeMux I__8595 (
            .O(N__40148),
            .I(N__40143));
    InMux I__8594 (
            .O(N__40147),
            .I(N__40140));
    InMux I__8593 (
            .O(N__40146),
            .I(N__40135));
    InMux I__8592 (
            .O(N__40143),
            .I(N__40135));
    LocalMux I__8591 (
            .O(N__40140),
            .I(N__40130));
    LocalMux I__8590 (
            .O(N__40135),
            .I(N__40130));
    Odrv4 I__8589 (
            .O(N__40130),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__8588 (
            .O(N__40127),
            .I(N__40124));
    LocalMux I__8587 (
            .O(N__40124),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    InMux I__8586 (
            .O(N__40121),
            .I(N__40118));
    LocalMux I__8585 (
            .O(N__40118),
            .I(N__40115));
    Span4Mux_v I__8584 (
            .O(N__40115),
            .I(N__40111));
    InMux I__8583 (
            .O(N__40114),
            .I(N__40108));
    Odrv4 I__8582 (
            .O(N__40111),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    LocalMux I__8581 (
            .O(N__40108),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__8580 (
            .O(N__40103),
            .I(N__40097));
    InMux I__8579 (
            .O(N__40102),
            .I(N__40097));
    LocalMux I__8578 (
            .O(N__40097),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    CascadeMux I__8577 (
            .O(N__40094),
            .I(N__40091));
    InMux I__8576 (
            .O(N__40091),
            .I(N__40088));
    LocalMux I__8575 (
            .O(N__40088),
            .I(N__40085));
    Odrv4 I__8574 (
            .O(N__40085),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    InMux I__8573 (
            .O(N__40082),
            .I(N__40079));
    LocalMux I__8572 (
            .O(N__40079),
            .I(N__40076));
    Span4Mux_h I__8571 (
            .O(N__40076),
            .I(N__40073));
    Odrv4 I__8570 (
            .O(N__40073),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    InMux I__8569 (
            .O(N__40070),
            .I(N__40064));
    InMux I__8568 (
            .O(N__40069),
            .I(N__40064));
    LocalMux I__8567 (
            .O(N__40064),
            .I(N__40060));
    InMux I__8566 (
            .O(N__40063),
            .I(N__40057));
    Span4Mux_h I__8565 (
            .O(N__40060),
            .I(N__40054));
    LocalMux I__8564 (
            .O(N__40057),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__8563 (
            .O(N__40054),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    CascadeMux I__8562 (
            .O(N__40049),
            .I(N__40046));
    InMux I__8561 (
            .O(N__40046),
            .I(N__40040));
    InMux I__8560 (
            .O(N__40045),
            .I(N__40040));
    LocalMux I__8559 (
            .O(N__40040),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    CascadeMux I__8558 (
            .O(N__40037),
            .I(N__40033));
    InMux I__8557 (
            .O(N__40036),
            .I(N__40028));
    InMux I__8556 (
            .O(N__40033),
            .I(N__40028));
    LocalMux I__8555 (
            .O(N__40028),
            .I(N__40024));
    InMux I__8554 (
            .O(N__40027),
            .I(N__40021));
    Span4Mux_h I__8553 (
            .O(N__40024),
            .I(N__40018));
    LocalMux I__8552 (
            .O(N__40021),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    Odrv4 I__8551 (
            .O(N__40018),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    CascadeMux I__8550 (
            .O(N__40013),
            .I(N__40010));
    InMux I__8549 (
            .O(N__40010),
            .I(N__40007));
    LocalMux I__8548 (
            .O(N__40007),
            .I(N__40004));
    Odrv4 I__8547 (
            .O(N__40004),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    InMux I__8546 (
            .O(N__40001),
            .I(N__39997));
    InMux I__8545 (
            .O(N__40000),
            .I(N__39993));
    LocalMux I__8544 (
            .O(N__39997),
            .I(N__39990));
    InMux I__8543 (
            .O(N__39996),
            .I(N__39987));
    LocalMux I__8542 (
            .O(N__39993),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv12 I__8541 (
            .O(N__39990),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    LocalMux I__8540 (
            .O(N__39987),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__8539 (
            .O(N__39980),
            .I(N__39974));
    InMux I__8538 (
            .O(N__39979),
            .I(N__39974));
    LocalMux I__8537 (
            .O(N__39974),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    InMux I__8536 (
            .O(N__39971),
            .I(N__39968));
    LocalMux I__8535 (
            .O(N__39968),
            .I(N__39964));
    InMux I__8534 (
            .O(N__39967),
            .I(N__39961));
    Odrv12 I__8533 (
            .O(N__39964),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__8532 (
            .O(N__39961),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    CascadeMux I__8531 (
            .O(N__39956),
            .I(N__39953));
    InMux I__8530 (
            .O(N__39953),
            .I(N__39950));
    LocalMux I__8529 (
            .O(N__39950),
            .I(N__39947));
    Odrv4 I__8528 (
            .O(N__39947),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    InMux I__8527 (
            .O(N__39944),
            .I(N__39938));
    InMux I__8526 (
            .O(N__39943),
            .I(N__39938));
    LocalMux I__8525 (
            .O(N__39938),
            .I(N__39934));
    InMux I__8524 (
            .O(N__39937),
            .I(N__39931));
    Span4Mux_h I__8523 (
            .O(N__39934),
            .I(N__39928));
    LocalMux I__8522 (
            .O(N__39931),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__8521 (
            .O(N__39928),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    CascadeMux I__8520 (
            .O(N__39923),
            .I(N__39920));
    InMux I__8519 (
            .O(N__39920),
            .I(N__39914));
    InMux I__8518 (
            .O(N__39919),
            .I(N__39914));
    LocalMux I__8517 (
            .O(N__39914),
            .I(N__39910));
    InMux I__8516 (
            .O(N__39913),
            .I(N__39907));
    Span4Mux_v I__8515 (
            .O(N__39910),
            .I(N__39904));
    LocalMux I__8514 (
            .O(N__39907),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__8513 (
            .O(N__39904),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__8512 (
            .O(N__39899),
            .I(N__39893));
    InMux I__8511 (
            .O(N__39898),
            .I(N__39893));
    LocalMux I__8510 (
            .O(N__39893),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    InMux I__8509 (
            .O(N__39890),
            .I(N__39887));
    LocalMux I__8508 (
            .O(N__39887),
            .I(N__39884));
    Span4Mux_h I__8507 (
            .O(N__39884),
            .I(N__39881));
    Odrv4 I__8506 (
            .O(N__39881),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    InMux I__8505 (
            .O(N__39878),
            .I(N__39875));
    LocalMux I__8504 (
            .O(N__39875),
            .I(N__39871));
    InMux I__8503 (
            .O(N__39874),
            .I(N__39868));
    Odrv12 I__8502 (
            .O(N__39871),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    LocalMux I__8501 (
            .O(N__39868),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    CascadeMux I__8500 (
            .O(N__39863),
            .I(N__39860));
    InMux I__8499 (
            .O(N__39860),
            .I(N__39854));
    InMux I__8498 (
            .O(N__39859),
            .I(N__39854));
    LocalMux I__8497 (
            .O(N__39854),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    CascadeMux I__8496 (
            .O(N__39851),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    CascadeMux I__8495 (
            .O(N__39848),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30_cascade_));
    InMux I__8494 (
            .O(N__39845),
            .I(N__39839));
    InMux I__8493 (
            .O(N__39844),
            .I(N__39839));
    LocalMux I__8492 (
            .O(N__39839),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    InMux I__8491 (
            .O(N__39836),
            .I(N__39831));
    InMux I__8490 (
            .O(N__39835),
            .I(N__39826));
    InMux I__8489 (
            .O(N__39834),
            .I(N__39826));
    LocalMux I__8488 (
            .O(N__39831),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__8487 (
            .O(N__39826),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__8486 (
            .O(N__39821),
            .I(N__39816));
    InMux I__8485 (
            .O(N__39820),
            .I(N__39811));
    InMux I__8484 (
            .O(N__39819),
            .I(N__39811));
    LocalMux I__8483 (
            .O(N__39816),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__8482 (
            .O(N__39811),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__8481 (
            .O(N__39806),
            .I(N__39803));
    LocalMux I__8480 (
            .O(N__39803),
            .I(N__39800));
    Span4Mux_h I__8479 (
            .O(N__39800),
            .I(N__39797));
    Odrv4 I__8478 (
            .O(N__39797),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    InMux I__8477 (
            .O(N__39794),
            .I(N__39791));
    LocalMux I__8476 (
            .O(N__39791),
            .I(N__39788));
    Span4Mux_h I__8475 (
            .O(N__39788),
            .I(N__39785));
    Odrv4 I__8474 (
            .O(N__39785),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__8473 (
            .O(N__39782),
            .I(N__39779));
    LocalMux I__8472 (
            .O(N__39779),
            .I(N__39776));
    Odrv4 I__8471 (
            .O(N__39776),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    InMux I__8470 (
            .O(N__39773),
            .I(N__39767));
    InMux I__8469 (
            .O(N__39772),
            .I(N__39767));
    LocalMux I__8468 (
            .O(N__39767),
            .I(N__39763));
    InMux I__8467 (
            .O(N__39766),
            .I(N__39760));
    Span4Mux_h I__8466 (
            .O(N__39763),
            .I(N__39757));
    LocalMux I__8465 (
            .O(N__39760),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__8464 (
            .O(N__39757),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__8463 (
            .O(N__39752),
            .I(N__39748));
    InMux I__8462 (
            .O(N__39751),
            .I(N__39743));
    InMux I__8461 (
            .O(N__39748),
            .I(N__39743));
    LocalMux I__8460 (
            .O(N__39743),
            .I(N__39739));
    InMux I__8459 (
            .O(N__39742),
            .I(N__39736));
    Span4Mux_h I__8458 (
            .O(N__39739),
            .I(N__39733));
    LocalMux I__8457 (
            .O(N__39736),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__8456 (
            .O(N__39733),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__8455 (
            .O(N__39728),
            .I(N__39725));
    InMux I__8454 (
            .O(N__39725),
            .I(N__39722));
    LocalMux I__8453 (
            .O(N__39722),
            .I(N__39719));
    Span4Mux_h I__8452 (
            .O(N__39719),
            .I(N__39716));
    Odrv4 I__8451 (
            .O(N__39716),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    InMux I__8450 (
            .O(N__39713),
            .I(N__39707));
    InMux I__8449 (
            .O(N__39712),
            .I(N__39707));
    LocalMux I__8448 (
            .O(N__39707),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__8447 (
            .O(N__39704),
            .I(N__39701));
    InMux I__8446 (
            .O(N__39701),
            .I(N__39695));
    InMux I__8445 (
            .O(N__39700),
            .I(N__39695));
    LocalMux I__8444 (
            .O(N__39695),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__8443 (
            .O(N__39692),
            .I(elapsed_time_ns_1_RNI69DN9_0_28_cascade_));
    InMux I__8442 (
            .O(N__39689),
            .I(N__39683));
    InMux I__8441 (
            .O(N__39688),
            .I(N__39683));
    LocalMux I__8440 (
            .O(N__39683),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    InMux I__8439 (
            .O(N__39680),
            .I(N__39677));
    LocalMux I__8438 (
            .O(N__39677),
            .I(N__39674));
    Span4Mux_v I__8437 (
            .O(N__39674),
            .I(N__39671));
    Odrv4 I__8436 (
            .O(N__39671),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    InMux I__8435 (
            .O(N__39668),
            .I(N__39663));
    InMux I__8434 (
            .O(N__39667),
            .I(N__39658));
    InMux I__8433 (
            .O(N__39666),
            .I(N__39658));
    LocalMux I__8432 (
            .O(N__39663),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__8431 (
            .O(N__39658),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    CascadeMux I__8430 (
            .O(N__39653),
            .I(N__39649));
    InMux I__8429 (
            .O(N__39652),
            .I(N__39645));
    InMux I__8428 (
            .O(N__39649),
            .I(N__39640));
    InMux I__8427 (
            .O(N__39648),
            .I(N__39640));
    LocalMux I__8426 (
            .O(N__39645),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__8425 (
            .O(N__39640),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    CascadeMux I__8424 (
            .O(N__39635),
            .I(N__39632));
    InMux I__8423 (
            .O(N__39632),
            .I(N__39629));
    LocalMux I__8422 (
            .O(N__39629),
            .I(N__39626));
    Span4Mux_v I__8421 (
            .O(N__39626),
            .I(N__39623));
    Span4Mux_h I__8420 (
            .O(N__39623),
            .I(N__39620));
    Odrv4 I__8419 (
            .O(N__39620),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    CascadeMux I__8418 (
            .O(N__39617),
            .I(elapsed_time_ns_1_RNI14DN9_0_23_cascade_));
    CascadeMux I__8417 (
            .O(N__39614),
            .I(N__39611));
    InMux I__8416 (
            .O(N__39611),
            .I(N__39605));
    InMux I__8415 (
            .O(N__39610),
            .I(N__39605));
    LocalMux I__8414 (
            .O(N__39605),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    CascadeMux I__8413 (
            .O(N__39602),
            .I(elapsed_time_ns_1_RNI03DN9_0_22_cascade_));
    InMux I__8412 (
            .O(N__39599),
            .I(N__39593));
    InMux I__8411 (
            .O(N__39598),
            .I(N__39593));
    LocalMux I__8410 (
            .O(N__39593),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    CascadeMux I__8409 (
            .O(N__39590),
            .I(N__39587));
    InMux I__8408 (
            .O(N__39587),
            .I(N__39584));
    LocalMux I__8407 (
            .O(N__39584),
            .I(N__39581));
    Span4Mux_h I__8406 (
            .O(N__39581),
            .I(N__39578));
    Odrv4 I__8405 (
            .O(N__39578),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__8404 (
            .O(N__39575),
            .I(N__39572));
    LocalMux I__8403 (
            .O(N__39572),
            .I(N__39568));
    InMux I__8402 (
            .O(N__39571),
            .I(N__39564));
    Span4Mux_v I__8401 (
            .O(N__39568),
            .I(N__39561));
    InMux I__8400 (
            .O(N__39567),
            .I(N__39558));
    LocalMux I__8399 (
            .O(N__39564),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__8398 (
            .O(N__39561),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    LocalMux I__8397 (
            .O(N__39558),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__8396 (
            .O(N__39551),
            .I(N__39546));
    InMux I__8395 (
            .O(N__39550),
            .I(N__39543));
    CascadeMux I__8394 (
            .O(N__39549),
            .I(N__39538));
    LocalMux I__8393 (
            .O(N__39546),
            .I(N__39535));
    LocalMux I__8392 (
            .O(N__39543),
            .I(N__39532));
    InMux I__8391 (
            .O(N__39542),
            .I(N__39527));
    InMux I__8390 (
            .O(N__39541),
            .I(N__39527));
    InMux I__8389 (
            .O(N__39538),
            .I(N__39524));
    Span4Mux_h I__8388 (
            .O(N__39535),
            .I(N__39521));
    Span4Mux_h I__8387 (
            .O(N__39532),
            .I(N__39518));
    LocalMux I__8386 (
            .O(N__39527),
            .I(N__39515));
    LocalMux I__8385 (
            .O(N__39524),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__8384 (
            .O(N__39521),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__8383 (
            .O(N__39518),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv12 I__8382 (
            .O(N__39515),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__8381 (
            .O(N__39506),
            .I(N__39501));
    InMux I__8380 (
            .O(N__39505),
            .I(N__39498));
    InMux I__8379 (
            .O(N__39504),
            .I(N__39495));
    LocalMux I__8378 (
            .O(N__39501),
            .I(N__39492));
    LocalMux I__8377 (
            .O(N__39498),
            .I(N__39489));
    LocalMux I__8376 (
            .O(N__39495),
            .I(N__39486));
    Span4Mux_h I__8375 (
            .O(N__39492),
            .I(N__39483));
    Odrv4 I__8374 (
            .O(N__39489),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__8373 (
            .O(N__39486),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__8372 (
            .O(N__39483),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__8371 (
            .O(N__39476),
            .I(N__39473));
    LocalMux I__8370 (
            .O(N__39473),
            .I(N__39470));
    Span4Mux_h I__8369 (
            .O(N__39470),
            .I(N__39466));
    InMux I__8368 (
            .O(N__39469),
            .I(N__39463));
    Odrv4 I__8367 (
            .O(N__39466),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__8366 (
            .O(N__39463),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__8365 (
            .O(N__39458),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__8364 (
            .O(N__39455),
            .I(N__39452));
    InMux I__8363 (
            .O(N__39452),
            .I(N__39447));
    InMux I__8362 (
            .O(N__39451),
            .I(N__39442));
    InMux I__8361 (
            .O(N__39450),
            .I(N__39442));
    LocalMux I__8360 (
            .O(N__39447),
            .I(N__39439));
    LocalMux I__8359 (
            .O(N__39442),
            .I(N__39434));
    Span4Mux_h I__8358 (
            .O(N__39439),
            .I(N__39431));
    InMux I__8357 (
            .O(N__39438),
            .I(N__39426));
    InMux I__8356 (
            .O(N__39437),
            .I(N__39426));
    Odrv4 I__8355 (
            .O(N__39434),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__8354 (
            .O(N__39431),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__8353 (
            .O(N__39426),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    InMux I__8352 (
            .O(N__39419),
            .I(N__39416));
    LocalMux I__8351 (
            .O(N__39416),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    CascadeMux I__8350 (
            .O(N__39413),
            .I(N__39410));
    InMux I__8349 (
            .O(N__39410),
            .I(N__39407));
    LocalMux I__8348 (
            .O(N__39407),
            .I(N__39404));
    Span4Mux_h I__8347 (
            .O(N__39404),
            .I(N__39401));
    Odrv4 I__8346 (
            .O(N__39401),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__8345 (
            .O(N__39398),
            .I(N__39391));
    InMux I__8344 (
            .O(N__39397),
            .I(N__39391));
    InMux I__8343 (
            .O(N__39396),
            .I(N__39388));
    LocalMux I__8342 (
            .O(N__39391),
            .I(N__39385));
    LocalMux I__8341 (
            .O(N__39388),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__8340 (
            .O(N__39385),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    CascadeMux I__8339 (
            .O(N__39380),
            .I(N__39377));
    InMux I__8338 (
            .O(N__39377),
            .I(N__39371));
    InMux I__8337 (
            .O(N__39376),
            .I(N__39371));
    LocalMux I__8336 (
            .O(N__39371),
            .I(N__39367));
    InMux I__8335 (
            .O(N__39370),
            .I(N__39364));
    Span4Mux_v I__8334 (
            .O(N__39367),
            .I(N__39361));
    LocalMux I__8333 (
            .O(N__39364),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__8332 (
            .O(N__39361),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__8331 (
            .O(N__39356),
            .I(N__39353));
    LocalMux I__8330 (
            .O(N__39353),
            .I(N__39350));
    Odrv4 I__8329 (
            .O(N__39350),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    CascadeMux I__8328 (
            .O(N__39347),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_));
    CascadeMux I__8327 (
            .O(N__39344),
            .I(N__39341));
    InMux I__8326 (
            .O(N__39341),
            .I(N__39335));
    InMux I__8325 (
            .O(N__39340),
            .I(N__39335));
    LocalMux I__8324 (
            .O(N__39335),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    InMux I__8323 (
            .O(N__39332),
            .I(N__39329));
    LocalMux I__8322 (
            .O(N__39329),
            .I(N__39326));
    Odrv4 I__8321 (
            .O(N__39326),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__8320 (
            .O(N__39323),
            .I(N__39320));
    LocalMux I__8319 (
            .O(N__39320),
            .I(N__39317));
    Odrv12 I__8318 (
            .O(N__39317),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    CascadeMux I__8317 (
            .O(N__39314),
            .I(N__39311));
    InMux I__8316 (
            .O(N__39311),
            .I(N__39308));
    LocalMux I__8315 (
            .O(N__39308),
            .I(N__39305));
    Span4Mux_v I__8314 (
            .O(N__39305),
            .I(N__39302));
    Odrv4 I__8313 (
            .O(N__39302),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__8312 (
            .O(N__39299),
            .I(N__39296));
    LocalMux I__8311 (
            .O(N__39296),
            .I(N__39293));
    Span4Mux_h I__8310 (
            .O(N__39293),
            .I(N__39289));
    InMux I__8309 (
            .O(N__39292),
            .I(N__39285));
    Span4Mux_v I__8308 (
            .O(N__39289),
            .I(N__39282));
    InMux I__8307 (
            .O(N__39288),
            .I(N__39279));
    LocalMux I__8306 (
            .O(N__39285),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    Odrv4 I__8305 (
            .O(N__39282),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    LocalMux I__8304 (
            .O(N__39279),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    InMux I__8303 (
            .O(N__39272),
            .I(N__39268));
    InMux I__8302 (
            .O(N__39271),
            .I(N__39265));
    LocalMux I__8301 (
            .O(N__39268),
            .I(N__39262));
    LocalMux I__8300 (
            .O(N__39265),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    Odrv4 I__8299 (
            .O(N__39262),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    CascadeMux I__8298 (
            .O(N__39257),
            .I(N__39252));
    InMux I__8297 (
            .O(N__39256),
            .I(N__39246));
    InMux I__8296 (
            .O(N__39255),
            .I(N__39246));
    InMux I__8295 (
            .O(N__39252),
            .I(N__39241));
    InMux I__8294 (
            .O(N__39251),
            .I(N__39241));
    LocalMux I__8293 (
            .O(N__39246),
            .I(N__39238));
    LocalMux I__8292 (
            .O(N__39241),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__8291 (
            .O(N__39238),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__8290 (
            .O(N__39233),
            .I(N__39229));
    InMux I__8289 (
            .O(N__39232),
            .I(N__39225));
    LocalMux I__8288 (
            .O(N__39229),
            .I(N__39222));
    InMux I__8287 (
            .O(N__39228),
            .I(N__39219));
    LocalMux I__8286 (
            .O(N__39225),
            .I(N__39214));
    Span4Mux_v I__8285 (
            .O(N__39222),
            .I(N__39214));
    LocalMux I__8284 (
            .O(N__39219),
            .I(N__39211));
    Odrv4 I__8283 (
            .O(N__39214),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv12 I__8282 (
            .O(N__39211),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    CascadeMux I__8281 (
            .O(N__39206),
            .I(N__39203));
    InMux I__8280 (
            .O(N__39203),
            .I(N__39200));
    LocalMux I__8279 (
            .O(N__39200),
            .I(N__39197));
    Odrv4 I__8278 (
            .O(N__39197),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ));
    CascadeMux I__8277 (
            .O(N__39194),
            .I(N__39191));
    InMux I__8276 (
            .O(N__39191),
            .I(N__39188));
    LocalMux I__8275 (
            .O(N__39188),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__8274 (
            .O(N__39185),
            .I(N__39182));
    LocalMux I__8273 (
            .O(N__39182),
            .I(N__39179));
    Odrv12 I__8272 (
            .O(N__39179),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    CascadeMux I__8271 (
            .O(N__39176),
            .I(N__39173));
    InMux I__8270 (
            .O(N__39173),
            .I(N__39170));
    LocalMux I__8269 (
            .O(N__39170),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__8268 (
            .O(N__39167),
            .I(N__39164));
    LocalMux I__8267 (
            .O(N__39164),
            .I(N__39161));
    Odrv4 I__8266 (
            .O(N__39161),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__8265 (
            .O(N__39158),
            .I(N__39155));
    LocalMux I__8264 (
            .O(N__39155),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__8263 (
            .O(N__39152),
            .I(N__39149));
    LocalMux I__8262 (
            .O(N__39149),
            .I(N__39146));
    Odrv4 I__8261 (
            .O(N__39146),
            .I(\current_shift_inst.control_input_axb_23 ));
    CascadeMux I__8260 (
            .O(N__39143),
            .I(N__39140));
    InMux I__8259 (
            .O(N__39140),
            .I(N__39137));
    LocalMux I__8258 (
            .O(N__39137),
            .I(N__39134));
    Odrv4 I__8257 (
            .O(N__39134),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    CascadeMux I__8256 (
            .O(N__39131),
            .I(N__39128));
    InMux I__8255 (
            .O(N__39128),
            .I(N__39125));
    LocalMux I__8254 (
            .O(N__39125),
            .I(N__39122));
    Span4Mux_v I__8253 (
            .O(N__39122),
            .I(N__39119));
    Odrv4 I__8252 (
            .O(N__39119),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    CascadeMux I__8251 (
            .O(N__39116),
            .I(N__39113));
    InMux I__8250 (
            .O(N__39113),
            .I(N__39110));
    LocalMux I__8249 (
            .O(N__39110),
            .I(N__39107));
    Span4Mux_h I__8248 (
            .O(N__39107),
            .I(N__39104));
    Odrv4 I__8247 (
            .O(N__39104),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    CascadeMux I__8246 (
            .O(N__39101),
            .I(N__39098));
    InMux I__8245 (
            .O(N__39098),
            .I(N__39095));
    LocalMux I__8244 (
            .O(N__39095),
            .I(N__39092));
    Odrv12 I__8243 (
            .O(N__39092),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    CascadeMux I__8242 (
            .O(N__39089),
            .I(N__39086));
    InMux I__8241 (
            .O(N__39086),
            .I(N__39083));
    LocalMux I__8240 (
            .O(N__39083),
            .I(N__39080));
    Span4Mux_v I__8239 (
            .O(N__39080),
            .I(N__39077));
    Odrv4 I__8238 (
            .O(N__39077),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    InMux I__8237 (
            .O(N__39074),
            .I(N__39071));
    LocalMux I__8236 (
            .O(N__39071),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__8235 (
            .O(N__39068),
            .I(N__39065));
    LocalMux I__8234 (
            .O(N__39065),
            .I(N__39062));
    Odrv12 I__8233 (
            .O(N__39062),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    InMux I__8232 (
            .O(N__39059),
            .I(N__39056));
    LocalMux I__8231 (
            .O(N__39056),
            .I(N__39053));
    Odrv4 I__8230 (
            .O(N__39053),
            .I(\current_shift_inst.control_input_axb_13 ));
    InMux I__8229 (
            .O(N__39050),
            .I(N__39047));
    LocalMux I__8228 (
            .O(N__39047),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__8227 (
            .O(N__39044),
            .I(N__39041));
    LocalMux I__8226 (
            .O(N__39041),
            .I(N__39038));
    Span4Mux_v I__8225 (
            .O(N__39038),
            .I(N__39035));
    Odrv4 I__8224 (
            .O(N__39035),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__8223 (
            .O(N__39032),
            .I(N__39029));
    LocalMux I__8222 (
            .O(N__39029),
            .I(N__39026));
    Odrv4 I__8221 (
            .O(N__39026),
            .I(\current_shift_inst.control_input_axb_14 ));
    InMux I__8220 (
            .O(N__39023),
            .I(N__39020));
    LocalMux I__8219 (
            .O(N__39020),
            .I(N__39017));
    Odrv4 I__8218 (
            .O(N__39017),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__8217 (
            .O(N__39014),
            .I(N__39011));
    LocalMux I__8216 (
            .O(N__39011),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__8215 (
            .O(N__39008),
            .I(N__39005));
    LocalMux I__8214 (
            .O(N__39005),
            .I(N__39002));
    Odrv4 I__8213 (
            .O(N__39002),
            .I(\current_shift_inst.control_input_axb_15 ));
    InMux I__8212 (
            .O(N__38999),
            .I(N__38996));
    LocalMux I__8211 (
            .O(N__38996),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__8210 (
            .O(N__38993),
            .I(N__38990));
    LocalMux I__8209 (
            .O(N__38990),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    CascadeMux I__8208 (
            .O(N__38987),
            .I(N__38984));
    InMux I__8207 (
            .O(N__38984),
            .I(N__38981));
    LocalMux I__8206 (
            .O(N__38981),
            .I(N__38978));
    Odrv12 I__8205 (
            .O(N__38978),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__8204 (
            .O(N__38975),
            .I(N__38972));
    LocalMux I__8203 (
            .O(N__38972),
            .I(N__38969));
    Odrv4 I__8202 (
            .O(N__38969),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    CascadeMux I__8201 (
            .O(N__38966),
            .I(N__38963));
    InMux I__8200 (
            .O(N__38963),
            .I(N__38960));
    LocalMux I__8199 (
            .O(N__38960),
            .I(N__38957));
    Odrv4 I__8198 (
            .O(N__38957),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__8197 (
            .O(N__38954),
            .I(N__38951));
    LocalMux I__8196 (
            .O(N__38951),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    CascadeMux I__8195 (
            .O(N__38948),
            .I(N__38945));
    InMux I__8194 (
            .O(N__38945),
            .I(N__38942));
    LocalMux I__8193 (
            .O(N__38942),
            .I(N__38939));
    Span4Mux_v I__8192 (
            .O(N__38939),
            .I(N__38936));
    Odrv4 I__8191 (
            .O(N__38936),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    CascadeMux I__8190 (
            .O(N__38933),
            .I(N__38930));
    InMux I__8189 (
            .O(N__38930),
            .I(N__38927));
    LocalMux I__8188 (
            .O(N__38927),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    CascadeMux I__8187 (
            .O(N__38924),
            .I(N__38921));
    InMux I__8186 (
            .O(N__38921),
            .I(N__38918));
    LocalMux I__8185 (
            .O(N__38918),
            .I(N__38915));
    Odrv4 I__8184 (
            .O(N__38915),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__8183 (
            .O(N__38912),
            .I(N__38909));
    LocalMux I__8182 (
            .O(N__38909),
            .I(N__38906));
    Odrv12 I__8181 (
            .O(N__38906),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__8180 (
            .O(N__38903),
            .I(N__38900));
    LocalMux I__8179 (
            .O(N__38900),
            .I(N__38897));
    Odrv4 I__8178 (
            .O(N__38897),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__8177 (
            .O(N__38894),
            .I(N__38891));
    LocalMux I__8176 (
            .O(N__38891),
            .I(N__38888));
    Odrv12 I__8175 (
            .O(N__38888),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__8174 (
            .O(N__38885),
            .I(N__38882));
    LocalMux I__8173 (
            .O(N__38882),
            .I(N__38879));
    Odrv12 I__8172 (
            .O(N__38879),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__8171 (
            .O(N__38876),
            .I(N__38873));
    LocalMux I__8170 (
            .O(N__38873),
            .I(N__38870));
    Odrv4 I__8169 (
            .O(N__38870),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__8168 (
            .O(N__38867),
            .I(N__38864));
    LocalMux I__8167 (
            .O(N__38864),
            .I(N__38861));
    Odrv12 I__8166 (
            .O(N__38861),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__8165 (
            .O(N__38858),
            .I(N__38855));
    LocalMux I__8164 (
            .O(N__38855),
            .I(N__38852));
    Odrv4 I__8163 (
            .O(N__38852),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__8162 (
            .O(N__38849),
            .I(N__38846));
    LocalMux I__8161 (
            .O(N__38846),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__8160 (
            .O(N__38843),
            .I(N__38840));
    LocalMux I__8159 (
            .O(N__38840),
            .I(N__38837));
    Span4Mux_v I__8158 (
            .O(N__38837),
            .I(N__38834));
    Odrv4 I__8157 (
            .O(N__38834),
            .I(\current_shift_inst.control_input_axb_24 ));
    InMux I__8156 (
            .O(N__38831),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__8155 (
            .O(N__38828),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__8154 (
            .O(N__38825),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__8153 (
            .O(N__38822),
            .I(N__38819));
    LocalMux I__8152 (
            .O(N__38819),
            .I(N__38816));
    Span4Mux_h I__8151 (
            .O(N__38816),
            .I(N__38813));
    Span4Mux_v I__8150 (
            .O(N__38813),
            .I(N__38810));
    Odrv4 I__8149 (
            .O(N__38810),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__8148 (
            .O(N__38807),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__8147 (
            .O(N__38804),
            .I(N__38801));
    LocalMux I__8146 (
            .O(N__38801),
            .I(N__38798));
    Span4Mux_v I__8145 (
            .O(N__38798),
            .I(N__38795));
    Sp12to4 I__8144 (
            .O(N__38795),
            .I(N__38792));
    Odrv12 I__8143 (
            .O(N__38792),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__8142 (
            .O(N__38789),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__8141 (
            .O(N__38786),
            .I(N__38783));
    LocalMux I__8140 (
            .O(N__38783),
            .I(N__38780));
    Span4Mux_h I__8139 (
            .O(N__38780),
            .I(N__38777));
    Odrv4 I__8138 (
            .O(N__38777),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__8137 (
            .O(N__38774),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__8136 (
            .O(N__38771),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__8135 (
            .O(N__38768),
            .I(N__38765));
    LocalMux I__8134 (
            .O(N__38765),
            .I(N__38762));
    Span4Mux_v I__8133 (
            .O(N__38762),
            .I(N__38759));
    Sp12to4 I__8132 (
            .O(N__38759),
            .I(N__38756));
    Odrv12 I__8131 (
            .O(N__38756),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__8130 (
            .O(N__38753),
            .I(N__38750));
    LocalMux I__8129 (
            .O(N__38750),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    InMux I__8128 (
            .O(N__38747),
            .I(N__38744));
    LocalMux I__8127 (
            .O(N__38744),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    InMux I__8126 (
            .O(N__38741),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    InMux I__8125 (
            .O(N__38738),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    CascadeMux I__8124 (
            .O(N__38735),
            .I(N__38732));
    InMux I__8123 (
            .O(N__38732),
            .I(N__38729));
    LocalMux I__8122 (
            .O(N__38729),
            .I(N__38726));
    Span4Mux_h I__8121 (
            .O(N__38726),
            .I(N__38723));
    Odrv4 I__8120 (
            .O(N__38723),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__8119 (
            .O(N__38720),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    CascadeMux I__8118 (
            .O(N__38717),
            .I(N__38714));
    InMux I__8117 (
            .O(N__38714),
            .I(N__38711));
    LocalMux I__8116 (
            .O(N__38711),
            .I(N__38708));
    Span4Mux_v I__8115 (
            .O(N__38708),
            .I(N__38705));
    Odrv4 I__8114 (
            .O(N__38705),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__8113 (
            .O(N__38702),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__8112 (
            .O(N__38699),
            .I(N__38696));
    LocalMux I__8111 (
            .O(N__38696),
            .I(N__38693));
    Span4Mux_v I__8110 (
            .O(N__38693),
            .I(N__38690));
    Odrv4 I__8109 (
            .O(N__38690),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__8108 (
            .O(N__38687),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__8107 (
            .O(N__38684),
            .I(N__38681));
    LocalMux I__8106 (
            .O(N__38681),
            .I(N__38678));
    Span4Mux_v I__8105 (
            .O(N__38678),
            .I(N__38675));
    Odrv4 I__8104 (
            .O(N__38675),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__8103 (
            .O(N__38672),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    CascadeMux I__8102 (
            .O(N__38669),
            .I(N__38666));
    InMux I__8101 (
            .O(N__38666),
            .I(N__38663));
    LocalMux I__8100 (
            .O(N__38663),
            .I(N__38660));
    Span4Mux_v I__8099 (
            .O(N__38660),
            .I(N__38657));
    Odrv4 I__8098 (
            .O(N__38657),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__8097 (
            .O(N__38654),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__8096 (
            .O(N__38651),
            .I(N__38648));
    LocalMux I__8095 (
            .O(N__38648),
            .I(N__38645));
    Span4Mux_v I__8094 (
            .O(N__38645),
            .I(N__38642));
    Odrv4 I__8093 (
            .O(N__38642),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__8092 (
            .O(N__38639),
            .I(bfn_15_16_0_));
    InMux I__8091 (
            .O(N__38636),
            .I(N__38633));
    LocalMux I__8090 (
            .O(N__38633),
            .I(N__38630));
    Span4Mux_v I__8089 (
            .O(N__38630),
            .I(N__38627));
    Odrv4 I__8088 (
            .O(N__38627),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__8087 (
            .O(N__38624),
            .I(N__38621));
    LocalMux I__8086 (
            .O(N__38621),
            .I(N__38618));
    Span4Mux_v I__8085 (
            .O(N__38618),
            .I(N__38615));
    Odrv4 I__8084 (
            .O(N__38615),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__8083 (
            .O(N__38612),
            .I(bfn_15_14_0_));
    InMux I__8082 (
            .O(N__38609),
            .I(N__38606));
    LocalMux I__8081 (
            .O(N__38606),
            .I(N__38603));
    Span4Mux_v I__8080 (
            .O(N__38603),
            .I(N__38600));
    Odrv4 I__8079 (
            .O(N__38600),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__8078 (
            .O(N__38597),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__8077 (
            .O(N__38594),
            .I(N__38591));
    LocalMux I__8076 (
            .O(N__38591),
            .I(N__38588));
    Span4Mux_v I__8075 (
            .O(N__38588),
            .I(N__38585));
    Odrv4 I__8074 (
            .O(N__38585),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__8073 (
            .O(N__38582),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__8072 (
            .O(N__38579),
            .I(N__38576));
    LocalMux I__8071 (
            .O(N__38576),
            .I(N__38573));
    Span4Mux_v I__8070 (
            .O(N__38573),
            .I(N__38570));
    Odrv4 I__8069 (
            .O(N__38570),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__8068 (
            .O(N__38567),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    InMux I__8067 (
            .O(N__38564),
            .I(N__38561));
    LocalMux I__8066 (
            .O(N__38561),
            .I(N__38558));
    Span12Mux_h I__8065 (
            .O(N__38558),
            .I(N__38555));
    Odrv12 I__8064 (
            .O(N__38555),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__8063 (
            .O(N__38552),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__8062 (
            .O(N__38549),
            .I(N__38546));
    LocalMux I__8061 (
            .O(N__38546),
            .I(N__38543));
    Span4Mux_v I__8060 (
            .O(N__38543),
            .I(N__38540));
    Odrv4 I__8059 (
            .O(N__38540),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__8058 (
            .O(N__38537),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    InMux I__8057 (
            .O(N__38534),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__8056 (
            .O(N__38531),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__8055 (
            .O(N__38528),
            .I(bfn_15_15_0_));
    CascadeMux I__8054 (
            .O(N__38525),
            .I(N__38522));
    InMux I__8053 (
            .O(N__38522),
            .I(N__38519));
    LocalMux I__8052 (
            .O(N__38519),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ));
    InMux I__8051 (
            .O(N__38516),
            .I(N__38513));
    LocalMux I__8050 (
            .O(N__38513),
            .I(N__38510));
    Span4Mux_v I__8049 (
            .O(N__38510),
            .I(N__38507));
    Span4Mux_h I__8048 (
            .O(N__38507),
            .I(N__38504));
    Odrv4 I__8047 (
            .O(N__38504),
            .I(\current_shift_inst.un38_control_input_0_s1_3 ));
    InMux I__8046 (
            .O(N__38501),
            .I(\current_shift_inst.un38_control_input_cry_2_s1 ));
    InMux I__8045 (
            .O(N__38498),
            .I(N__38495));
    LocalMux I__8044 (
            .O(N__38495),
            .I(N__38492));
    Span4Mux_v I__8043 (
            .O(N__38492),
            .I(N__38489));
    Span4Mux_v I__8042 (
            .O(N__38489),
            .I(N__38486));
    Odrv4 I__8041 (
            .O(N__38486),
            .I(\current_shift_inst.un38_control_input_0_s1_4 ));
    InMux I__8040 (
            .O(N__38483),
            .I(\current_shift_inst.un38_control_input_cry_3_s1 ));
    CascadeMux I__8039 (
            .O(N__38480),
            .I(N__38477));
    InMux I__8038 (
            .O(N__38477),
            .I(N__38474));
    LocalMux I__8037 (
            .O(N__38474),
            .I(N__38471));
    Span12Mux_h I__8036 (
            .O(N__38471),
            .I(N__38468));
    Odrv12 I__8035 (
            .O(N__38468),
            .I(\current_shift_inst.un38_control_input_0_s1_5 ));
    InMux I__8034 (
            .O(N__38465),
            .I(\current_shift_inst.un38_control_input_cry_4_s1 ));
    InMux I__8033 (
            .O(N__38462),
            .I(N__38459));
    LocalMux I__8032 (
            .O(N__38459),
            .I(N__38456));
    Span12Mux_v I__8031 (
            .O(N__38456),
            .I(N__38453));
    Odrv12 I__8030 (
            .O(N__38453),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__8029 (
            .O(N__38450),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__8028 (
            .O(N__38447),
            .I(N__38444));
    LocalMux I__8027 (
            .O(N__38444),
            .I(N__38441));
    Span4Mux_h I__8026 (
            .O(N__38441),
            .I(N__38438));
    Span4Mux_v I__8025 (
            .O(N__38438),
            .I(N__38435));
    Odrv4 I__8024 (
            .O(N__38435),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__8023 (
            .O(N__38432),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    InMux I__8022 (
            .O(N__38429),
            .I(N__38426));
    LocalMux I__8021 (
            .O(N__38426),
            .I(N__38423));
    Span4Mux_v I__8020 (
            .O(N__38423),
            .I(N__38420));
    Odrv4 I__8019 (
            .O(N__38420),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    CascadeMux I__8018 (
            .O(N__38417),
            .I(N__38414));
    InMux I__8017 (
            .O(N__38414),
            .I(N__38411));
    LocalMux I__8016 (
            .O(N__38411),
            .I(N__38408));
    Span4Mux_v I__8015 (
            .O(N__38408),
            .I(N__38405));
    Odrv4 I__8014 (
            .O(N__38405),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    InMux I__8013 (
            .O(N__38402),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    CascadeMux I__8012 (
            .O(N__38399),
            .I(N__38396));
    InMux I__8011 (
            .O(N__38396),
            .I(N__38393));
    LocalMux I__8010 (
            .O(N__38393),
            .I(N__38388));
    InMux I__8009 (
            .O(N__38392),
            .I(N__38385));
    InMux I__8008 (
            .O(N__38391),
            .I(N__38382));
    Span4Mux_h I__8007 (
            .O(N__38388),
            .I(N__38379));
    LocalMux I__8006 (
            .O(N__38385),
            .I(N__38376));
    LocalMux I__8005 (
            .O(N__38382),
            .I(N__38373));
    Span4Mux_h I__8004 (
            .O(N__38379),
            .I(N__38370));
    Span4Mux_h I__8003 (
            .O(N__38376),
            .I(N__38367));
    Span4Mux_v I__8002 (
            .O(N__38373),
            .I(N__38364));
    Span4Mux_v I__8001 (
            .O(N__38370),
            .I(N__38361));
    Span4Mux_h I__8000 (
            .O(N__38367),
            .I(N__38358));
    Odrv4 I__7999 (
            .O(N__38364),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__7998 (
            .O(N__38361),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__7997 (
            .O(N__38358),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__7996 (
            .O(N__38351),
            .I(N__38348));
    LocalMux I__7995 (
            .O(N__38348),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    InMux I__7994 (
            .O(N__38345),
            .I(N__38341));
    InMux I__7993 (
            .O(N__38344),
            .I(N__38338));
    LocalMux I__7992 (
            .O(N__38341),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__7991 (
            .O(N__38338),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__7990 (
            .O(N__38333),
            .I(N__38330));
    InMux I__7989 (
            .O(N__38330),
            .I(N__38327));
    LocalMux I__7988 (
            .O(N__38327),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__7987 (
            .O(N__38324),
            .I(N__38320));
    InMux I__7986 (
            .O(N__38323),
            .I(N__38317));
    LocalMux I__7985 (
            .O(N__38320),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__7984 (
            .O(N__38317),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__7983 (
            .O(N__38312),
            .I(N__38309));
    InMux I__7982 (
            .O(N__38309),
            .I(N__38306));
    LocalMux I__7981 (
            .O(N__38306),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__7980 (
            .O(N__38303),
            .I(N__38299));
    InMux I__7979 (
            .O(N__38302),
            .I(N__38296));
    LocalMux I__7978 (
            .O(N__38299),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__7977 (
            .O(N__38296),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__7976 (
            .O(N__38291),
            .I(N__38288));
    InMux I__7975 (
            .O(N__38288),
            .I(N__38285));
    LocalMux I__7974 (
            .O(N__38285),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__7973 (
            .O(N__38282),
            .I(N__38278));
    InMux I__7972 (
            .O(N__38281),
            .I(N__38275));
    LocalMux I__7971 (
            .O(N__38278),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__7970 (
            .O(N__38275),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__7969 (
            .O(N__38270),
            .I(N__38267));
    InMux I__7968 (
            .O(N__38267),
            .I(N__38264));
    LocalMux I__7967 (
            .O(N__38264),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__7966 (
            .O(N__38261),
            .I(N__38257));
    InMux I__7965 (
            .O(N__38260),
            .I(N__38254));
    LocalMux I__7964 (
            .O(N__38257),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__7963 (
            .O(N__38254),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__7962 (
            .O(N__38249),
            .I(N__38246));
    InMux I__7961 (
            .O(N__38246),
            .I(N__38243));
    LocalMux I__7960 (
            .O(N__38243),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__7959 (
            .O(N__38240),
            .I(N__38236));
    InMux I__7958 (
            .O(N__38239),
            .I(N__38233));
    LocalMux I__7957 (
            .O(N__38236),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__7956 (
            .O(N__38233),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__7955 (
            .O(N__38228),
            .I(N__38225));
    InMux I__7954 (
            .O(N__38225),
            .I(N__38222));
    LocalMux I__7953 (
            .O(N__38222),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__7952 (
            .O(N__38219),
            .I(N__38215));
    InMux I__7951 (
            .O(N__38218),
            .I(N__38212));
    LocalMux I__7950 (
            .O(N__38215),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__7949 (
            .O(N__38212),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__7948 (
            .O(N__38207),
            .I(N__38204));
    LocalMux I__7947 (
            .O(N__38204),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__7946 (
            .O(N__38201),
            .I(N__38198));
    InMux I__7945 (
            .O(N__38198),
            .I(N__38195));
    LocalMux I__7944 (
            .O(N__38195),
            .I(N__38192));
    Odrv4 I__7943 (
            .O(N__38192),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    InMux I__7942 (
            .O(N__38189),
            .I(N__38185));
    InMux I__7941 (
            .O(N__38188),
            .I(N__38182));
    LocalMux I__7940 (
            .O(N__38185),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__7939 (
            .O(N__38182),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__7938 (
            .O(N__38177),
            .I(N__38174));
    LocalMux I__7937 (
            .O(N__38174),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__7936 (
            .O(N__38171),
            .I(N__38168));
    InMux I__7935 (
            .O(N__38168),
            .I(N__38165));
    LocalMux I__7934 (
            .O(N__38165),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__7933 (
            .O(N__38162),
            .I(N__38158));
    InMux I__7932 (
            .O(N__38161),
            .I(N__38154));
    InMux I__7931 (
            .O(N__38158),
            .I(N__38151));
    InMux I__7930 (
            .O(N__38157),
            .I(N__38148));
    LocalMux I__7929 (
            .O(N__38154),
            .I(N__38145));
    LocalMux I__7928 (
            .O(N__38151),
            .I(N__38142));
    LocalMux I__7927 (
            .O(N__38148),
            .I(N__38137));
    Span4Mux_h I__7926 (
            .O(N__38145),
            .I(N__38137));
    Odrv12 I__7925 (
            .O(N__38142),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__7924 (
            .O(N__38137),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__7923 (
            .O(N__38132),
            .I(N__38129));
    LocalMux I__7922 (
            .O(N__38129),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__7921 (
            .O(N__38126),
            .I(N__38123));
    LocalMux I__7920 (
            .O(N__38123),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    InMux I__7919 (
            .O(N__38120),
            .I(N__38116));
    InMux I__7918 (
            .O(N__38119),
            .I(N__38113));
    LocalMux I__7917 (
            .O(N__38116),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__7916 (
            .O(N__38113),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__7915 (
            .O(N__38108),
            .I(N__38105));
    InMux I__7914 (
            .O(N__38105),
            .I(N__38102));
    LocalMux I__7913 (
            .O(N__38102),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__7912 (
            .O(N__38099),
            .I(N__38096));
    InMux I__7911 (
            .O(N__38096),
            .I(N__38093));
    LocalMux I__7910 (
            .O(N__38093),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    InMux I__7909 (
            .O(N__38090),
            .I(N__38086));
    InMux I__7908 (
            .O(N__38089),
            .I(N__38083));
    LocalMux I__7907 (
            .O(N__38086),
            .I(N__38080));
    LocalMux I__7906 (
            .O(N__38083),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__7905 (
            .O(N__38080),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__7904 (
            .O(N__38075),
            .I(N__38072));
    LocalMux I__7903 (
            .O(N__38072),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__7902 (
            .O(N__38069),
            .I(N__38065));
    InMux I__7901 (
            .O(N__38068),
            .I(N__38062));
    LocalMux I__7900 (
            .O(N__38065),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__7899 (
            .O(N__38062),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__7898 (
            .O(N__38057),
            .I(N__38054));
    LocalMux I__7897 (
            .O(N__38054),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__7896 (
            .O(N__38051),
            .I(N__38048));
    InMux I__7895 (
            .O(N__38048),
            .I(N__38045));
    LocalMux I__7894 (
            .O(N__38045),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__7893 (
            .O(N__38042),
            .I(N__38039));
    LocalMux I__7892 (
            .O(N__38039),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    InMux I__7891 (
            .O(N__38036),
            .I(N__38032));
    InMux I__7890 (
            .O(N__38035),
            .I(N__38029));
    LocalMux I__7889 (
            .O(N__38032),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__7888 (
            .O(N__38029),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__7887 (
            .O(N__38024),
            .I(N__38021));
    InMux I__7886 (
            .O(N__38021),
            .I(N__38018));
    LocalMux I__7885 (
            .O(N__38018),
            .I(N__38015));
    Odrv4 I__7884 (
            .O(N__38015),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__7883 (
            .O(N__38012),
            .I(N__38008));
    InMux I__7882 (
            .O(N__38011),
            .I(N__38005));
    LocalMux I__7881 (
            .O(N__38008),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__7880 (
            .O(N__38005),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__7879 (
            .O(N__38000),
            .I(N__37997));
    LocalMux I__7878 (
            .O(N__37997),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__7877 (
            .O(N__37994),
            .I(N__37991));
    InMux I__7876 (
            .O(N__37991),
            .I(N__37988));
    LocalMux I__7875 (
            .O(N__37988),
            .I(N__37985));
    Odrv4 I__7874 (
            .O(N__37985),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__7873 (
            .O(N__37982),
            .I(N__37978));
    InMux I__7872 (
            .O(N__37981),
            .I(N__37975));
    LocalMux I__7871 (
            .O(N__37978),
            .I(N__37972));
    LocalMux I__7870 (
            .O(N__37975),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__7869 (
            .O(N__37972),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__7868 (
            .O(N__37967),
            .I(N__37964));
    LocalMux I__7867 (
            .O(N__37964),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__7866 (
            .O(N__37961),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__7865 (
            .O(N__37958),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__7864 (
            .O(N__37955),
            .I(N__37952));
    LocalMux I__7863 (
            .O(N__37952),
            .I(N__37949));
    Span4Mux_h I__7862 (
            .O(N__37949),
            .I(N__37945));
    InMux I__7861 (
            .O(N__37948),
            .I(N__37942));
    Odrv4 I__7860 (
            .O(N__37945),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__7859 (
            .O(N__37942),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    InMux I__7858 (
            .O(N__37937),
            .I(N__37932));
    InMux I__7857 (
            .O(N__37936),
            .I(N__37929));
    InMux I__7856 (
            .O(N__37935),
            .I(N__37926));
    LocalMux I__7855 (
            .O(N__37932),
            .I(N__37923));
    LocalMux I__7854 (
            .O(N__37929),
            .I(N__37918));
    LocalMux I__7853 (
            .O(N__37926),
            .I(N__37918));
    Odrv12 I__7852 (
            .O(N__37923),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    Odrv4 I__7851 (
            .O(N__37918),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    InMux I__7850 (
            .O(N__37913),
            .I(N__37908));
    InMux I__7849 (
            .O(N__37912),
            .I(N__37905));
    InMux I__7848 (
            .O(N__37911),
            .I(N__37902));
    LocalMux I__7847 (
            .O(N__37908),
            .I(N__37899));
    LocalMux I__7846 (
            .O(N__37905),
            .I(N__37896));
    LocalMux I__7845 (
            .O(N__37902),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv4 I__7844 (
            .O(N__37899),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv4 I__7843 (
            .O(N__37896),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    InMux I__7842 (
            .O(N__37889),
            .I(N__37885));
    InMux I__7841 (
            .O(N__37888),
            .I(N__37882));
    LocalMux I__7840 (
            .O(N__37885),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__7839 (
            .O(N__37882),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__7838 (
            .O(N__37877),
            .I(N__37873));
    InMux I__7837 (
            .O(N__37876),
            .I(N__37869));
    LocalMux I__7836 (
            .O(N__37873),
            .I(N__37866));
    InMux I__7835 (
            .O(N__37872),
            .I(N__37863));
    LocalMux I__7834 (
            .O(N__37869),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__7833 (
            .O(N__37866),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    LocalMux I__7832 (
            .O(N__37863),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    InMux I__7831 (
            .O(N__37856),
            .I(N__37852));
    InMux I__7830 (
            .O(N__37855),
            .I(N__37848));
    LocalMux I__7829 (
            .O(N__37852),
            .I(N__37845));
    InMux I__7828 (
            .O(N__37851),
            .I(N__37842));
    LocalMux I__7827 (
            .O(N__37848),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__7826 (
            .O(N__37845),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__7825 (
            .O(N__37842),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__7824 (
            .O(N__37835),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__7823 (
            .O(N__37832),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__7822 (
            .O(N__37829),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__7821 (
            .O(N__37826),
            .I(N__37823));
    LocalMux I__7820 (
            .O(N__37823),
            .I(N__37818));
    InMux I__7819 (
            .O(N__37822),
            .I(N__37815));
    InMux I__7818 (
            .O(N__37821),
            .I(N__37812));
    Span4Mux_h I__7817 (
            .O(N__37818),
            .I(N__37809));
    LocalMux I__7816 (
            .O(N__37815),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__7815 (
            .O(N__37812),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__7814 (
            .O(N__37809),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__7813 (
            .O(N__37802),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__7812 (
            .O(N__37799),
            .I(N__37795));
    CascadeMux I__7811 (
            .O(N__37798),
            .I(N__37791));
    LocalMux I__7810 (
            .O(N__37795),
            .I(N__37788));
    InMux I__7809 (
            .O(N__37794),
            .I(N__37785));
    InMux I__7808 (
            .O(N__37791),
            .I(N__37782));
    Span4Mux_h I__7807 (
            .O(N__37788),
            .I(N__37779));
    LocalMux I__7806 (
            .O(N__37785),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__7805 (
            .O(N__37782),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__7804 (
            .O(N__37779),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__7803 (
            .O(N__37772),
            .I(bfn_15_8_0_));
    CascadeMux I__7802 (
            .O(N__37769),
            .I(N__37765));
    InMux I__7801 (
            .O(N__37768),
            .I(N__37761));
    InMux I__7800 (
            .O(N__37765),
            .I(N__37756));
    InMux I__7799 (
            .O(N__37764),
            .I(N__37756));
    LocalMux I__7798 (
            .O(N__37761),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__7797 (
            .O(N__37756),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__7796 (
            .O(N__37751),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__7795 (
            .O(N__37748),
            .I(N__37743));
    InMux I__7794 (
            .O(N__37747),
            .I(N__37738));
    InMux I__7793 (
            .O(N__37746),
            .I(N__37738));
    LocalMux I__7792 (
            .O(N__37743),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__7791 (
            .O(N__37738),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__7790 (
            .O(N__37733),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__7789 (
            .O(N__37730),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__7788 (
            .O(N__37727),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__7787 (
            .O(N__37724),
            .I(N__37720));
    InMux I__7786 (
            .O(N__37723),
            .I(N__37717));
    LocalMux I__7785 (
            .O(N__37720),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__7784 (
            .O(N__37717),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__7783 (
            .O(N__37712),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__7782 (
            .O(N__37709),
            .I(N__37705));
    InMux I__7781 (
            .O(N__37708),
            .I(N__37702));
    LocalMux I__7780 (
            .O(N__37705),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__7779 (
            .O(N__37702),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__7778 (
            .O(N__37697),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__7777 (
            .O(N__37694),
            .I(N__37690));
    InMux I__7776 (
            .O(N__37693),
            .I(N__37687));
    LocalMux I__7775 (
            .O(N__37690),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__7774 (
            .O(N__37687),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__7773 (
            .O(N__37682),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__7772 (
            .O(N__37679),
            .I(N__37675));
    InMux I__7771 (
            .O(N__37678),
            .I(N__37672));
    LocalMux I__7770 (
            .O(N__37675),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__7769 (
            .O(N__37672),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__7768 (
            .O(N__37667),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__7767 (
            .O(N__37664),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__7766 (
            .O(N__37661),
            .I(bfn_15_7_0_));
    CascadeMux I__7765 (
            .O(N__37658),
            .I(N__37654));
    InMux I__7764 (
            .O(N__37657),
            .I(N__37650));
    InMux I__7763 (
            .O(N__37654),
            .I(N__37647));
    InMux I__7762 (
            .O(N__37653),
            .I(N__37644));
    LocalMux I__7761 (
            .O(N__37650),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__7760 (
            .O(N__37647),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__7759 (
            .O(N__37644),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__7758 (
            .O(N__37637),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__7757 (
            .O(N__37634),
            .I(N__37629));
    InMux I__7756 (
            .O(N__37633),
            .I(N__37626));
    InMux I__7755 (
            .O(N__37632),
            .I(N__37623));
    LocalMux I__7754 (
            .O(N__37629),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__7753 (
            .O(N__37626),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__7752 (
            .O(N__37623),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__7751 (
            .O(N__37616),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    CascadeMux I__7750 (
            .O(N__37613),
            .I(N__37609));
    CascadeMux I__7749 (
            .O(N__37612),
            .I(N__37605));
    InMux I__7748 (
            .O(N__37609),
            .I(N__37602));
    InMux I__7747 (
            .O(N__37608),
            .I(N__37599));
    InMux I__7746 (
            .O(N__37605),
            .I(N__37596));
    LocalMux I__7745 (
            .O(N__37602),
            .I(N__37593));
    LocalMux I__7744 (
            .O(N__37599),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    LocalMux I__7743 (
            .O(N__37596),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__7742 (
            .O(N__37593),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__7741 (
            .O(N__37586),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__7740 (
            .O(N__37583),
            .I(N__37579));
    InMux I__7739 (
            .O(N__37582),
            .I(N__37576));
    LocalMux I__7738 (
            .O(N__37579),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__7737 (
            .O(N__37576),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__7736 (
            .O(N__37571),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__7735 (
            .O(N__37568),
            .I(N__37564));
    InMux I__7734 (
            .O(N__37567),
            .I(N__37561));
    LocalMux I__7733 (
            .O(N__37564),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__7732 (
            .O(N__37561),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__7731 (
            .O(N__37556),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__7730 (
            .O(N__37553),
            .I(N__37549));
    InMux I__7729 (
            .O(N__37552),
            .I(N__37546));
    LocalMux I__7728 (
            .O(N__37549),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__7727 (
            .O(N__37546),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__7726 (
            .O(N__37541),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__7725 (
            .O(N__37538),
            .I(N__37534));
    InMux I__7724 (
            .O(N__37537),
            .I(N__37531));
    LocalMux I__7723 (
            .O(N__37534),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__7722 (
            .O(N__37531),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__7721 (
            .O(N__37526),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__7720 (
            .O(N__37523),
            .I(N__37519));
    InMux I__7719 (
            .O(N__37522),
            .I(N__37516));
    LocalMux I__7718 (
            .O(N__37519),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__7717 (
            .O(N__37516),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__7716 (
            .O(N__37511),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__7715 (
            .O(N__37508),
            .I(N__37504));
    InMux I__7714 (
            .O(N__37507),
            .I(N__37501));
    LocalMux I__7713 (
            .O(N__37504),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__7712 (
            .O(N__37501),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__7711 (
            .O(N__37496),
            .I(bfn_15_6_0_));
    InMux I__7710 (
            .O(N__37493),
            .I(N__37489));
    InMux I__7709 (
            .O(N__37492),
            .I(N__37486));
    LocalMux I__7708 (
            .O(N__37489),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__7707 (
            .O(N__37486),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__7706 (
            .O(N__37481),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__7705 (
            .O(N__37478),
            .I(N__37474));
    InMux I__7704 (
            .O(N__37477),
            .I(N__37471));
    LocalMux I__7703 (
            .O(N__37474),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__7702 (
            .O(N__37471),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__7701 (
            .O(N__37466),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__7700 (
            .O(N__37463),
            .I(N__37457));
    InMux I__7699 (
            .O(N__37462),
            .I(N__37452));
    InMux I__7698 (
            .O(N__37461),
            .I(N__37452));
    InMux I__7697 (
            .O(N__37460),
            .I(N__37449));
    LocalMux I__7696 (
            .O(N__37457),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7695 (
            .O(N__37452),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7694 (
            .O(N__37449),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__7693 (
            .O(N__37442),
            .I(N__37436));
    InMux I__7692 (
            .O(N__37441),
            .I(N__37431));
    InMux I__7691 (
            .O(N__37440),
            .I(N__37431));
    InMux I__7690 (
            .O(N__37439),
            .I(N__37428));
    LocalMux I__7689 (
            .O(N__37436),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7688 (
            .O(N__37431),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7687 (
            .O(N__37428),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    CascadeMux I__7686 (
            .O(N__37421),
            .I(N__37417));
    InMux I__7685 (
            .O(N__37420),
            .I(N__37412));
    InMux I__7684 (
            .O(N__37417),
            .I(N__37409));
    InMux I__7683 (
            .O(N__37416),
            .I(N__37406));
    InMux I__7682 (
            .O(N__37415),
            .I(N__37403));
    LocalMux I__7681 (
            .O(N__37412),
            .I(N__37400));
    LocalMux I__7680 (
            .O(N__37409),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7679 (
            .O(N__37406),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7678 (
            .O(N__37403),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__7677 (
            .O(N__37400),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    CascadeMux I__7676 (
            .O(N__37391),
            .I(N__37388));
    InMux I__7675 (
            .O(N__37388),
            .I(N__37385));
    LocalMux I__7674 (
            .O(N__37385),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__7673 (
            .O(N__37382),
            .I(N__37379));
    LocalMux I__7672 (
            .O(N__37379),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__7671 (
            .O(N__37376),
            .I(N__37373));
    LocalMux I__7670 (
            .O(N__37373),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__7669 (
            .O(N__37370),
            .I(N__37367));
    LocalMux I__7668 (
            .O(N__37367),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__7667 (
            .O(N__37364),
            .I(N__37360));
    InMux I__7666 (
            .O(N__37363),
            .I(N__37355));
    InMux I__7665 (
            .O(N__37360),
            .I(N__37355));
    LocalMux I__7664 (
            .O(N__37355),
            .I(N__37352));
    Odrv4 I__7663 (
            .O(N__37352),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    CascadeMux I__7662 (
            .O(N__37349),
            .I(N__37346));
    InMux I__7661 (
            .O(N__37346),
            .I(N__37342));
    CascadeMux I__7660 (
            .O(N__37345),
            .I(N__37339));
    LocalMux I__7659 (
            .O(N__37342),
            .I(N__37336));
    InMux I__7658 (
            .O(N__37339),
            .I(N__37332));
    Span4Mux_v I__7657 (
            .O(N__37336),
            .I(N__37329));
    InMux I__7656 (
            .O(N__37335),
            .I(N__37326));
    LocalMux I__7655 (
            .O(N__37332),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__7654 (
            .O(N__37329),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__7653 (
            .O(N__37326),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__7652 (
            .O(N__37319),
            .I(N__37315));
    InMux I__7651 (
            .O(N__37318),
            .I(N__37312));
    LocalMux I__7650 (
            .O(N__37315),
            .I(N__37309));
    LocalMux I__7649 (
            .O(N__37312),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__7648 (
            .O(N__37309),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__7647 (
            .O(N__37304),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__7646 (
            .O(N__37301),
            .I(N__37297));
    InMux I__7645 (
            .O(N__37300),
            .I(N__37294));
    LocalMux I__7644 (
            .O(N__37297),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__7643 (
            .O(N__37294),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__7642 (
            .O(N__37289),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    CascadeMux I__7641 (
            .O(N__37286),
            .I(N__37283));
    InMux I__7640 (
            .O(N__37283),
            .I(N__37280));
    LocalMux I__7639 (
            .O(N__37280),
            .I(N__37277));
    Odrv4 I__7638 (
            .O(N__37277),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    CascadeMux I__7637 (
            .O(N__37274),
            .I(N__37271));
    InMux I__7636 (
            .O(N__37271),
            .I(N__37268));
    LocalMux I__7635 (
            .O(N__37268),
            .I(N__37265));
    Odrv4 I__7634 (
            .O(N__37265),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    CascadeMux I__7633 (
            .O(N__37262),
            .I(N__37259));
    InMux I__7632 (
            .O(N__37259),
            .I(N__37256));
    LocalMux I__7631 (
            .O(N__37256),
            .I(N__37253));
    Odrv4 I__7630 (
            .O(N__37253),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    InMux I__7629 (
            .O(N__37250),
            .I(N__37247));
    LocalMux I__7628 (
            .O(N__37247),
            .I(N__37244));
    Odrv4 I__7627 (
            .O(N__37244),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__7626 (
            .O(N__37241),
            .I(N__37238));
    LocalMux I__7625 (
            .O(N__37238),
            .I(N__37235));
    Odrv4 I__7624 (
            .O(N__37235),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__7623 (
            .O(N__37232),
            .I(N__37229));
    LocalMux I__7622 (
            .O(N__37229),
            .I(N__37226));
    Odrv4 I__7621 (
            .O(N__37226),
            .I(\current_shift_inst.control_input_axb_19 ));
    InMux I__7620 (
            .O(N__37223),
            .I(N__37220));
    LocalMux I__7619 (
            .O(N__37220),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__7618 (
            .O(N__37217),
            .I(N__37214));
    LocalMux I__7617 (
            .O(N__37214),
            .I(N__37211));
    Odrv12 I__7616 (
            .O(N__37211),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__7615 (
            .O(N__37208),
            .I(N__37205));
    LocalMux I__7614 (
            .O(N__37205),
            .I(N__37202));
    Odrv4 I__7613 (
            .O(N__37202),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__7612 (
            .O(N__37199),
            .I(N__37196));
    LocalMux I__7611 (
            .O(N__37196),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__7610 (
            .O(N__37193),
            .I(bfn_14_18_0_));
    InMux I__7609 (
            .O(N__37190),
            .I(N__37187));
    LocalMux I__7608 (
            .O(N__37187),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__7607 (
            .O(N__37184),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__7606 (
            .O(N__37181),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__7605 (
            .O(N__37178),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__7604 (
            .O(N__37175),
            .I(N__37172));
    LocalMux I__7603 (
            .O(N__37172),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__7602 (
            .O(N__37169),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__7601 (
            .O(N__37166),
            .I(N__37163));
    LocalMux I__7600 (
            .O(N__37163),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__7599 (
            .O(N__37160),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__7598 (
            .O(N__37157),
            .I(N__37154));
    LocalMux I__7597 (
            .O(N__37154),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__7596 (
            .O(N__37151),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__7595 (
            .O(N__37148),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__7594 (
            .O(N__37145),
            .I(N__37142));
    LocalMux I__7593 (
            .O(N__37142),
            .I(N__37139));
    Span4Mux_h I__7592 (
            .O(N__37139),
            .I(N__37136));
    Odrv4 I__7591 (
            .O(N__37136),
            .I(\current_shift_inst.control_input_axb_28 ));
    InMux I__7590 (
            .O(N__37133),
            .I(N__37130));
    LocalMux I__7589 (
            .O(N__37130),
            .I(N__37127));
    Odrv12 I__7588 (
            .O(N__37127),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    InMux I__7587 (
            .O(N__37124),
            .I(bfn_14_17_0_));
    InMux I__7586 (
            .O(N__37121),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    InMux I__7585 (
            .O(N__37118),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__7584 (
            .O(N__37115),
            .I(N__37112));
    LocalMux I__7583 (
            .O(N__37112),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__7582 (
            .O(N__37109),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    InMux I__7581 (
            .O(N__37106),
            .I(N__37103));
    LocalMux I__7580 (
            .O(N__37103),
            .I(N__37100));
    Odrv4 I__7579 (
            .O(N__37100),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__7578 (
            .O(N__37097),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__7577 (
            .O(N__37094),
            .I(N__37091));
    LocalMux I__7576 (
            .O(N__37091),
            .I(N__37088));
    Sp12to4 I__7575 (
            .O(N__37088),
            .I(N__37085));
    Odrv12 I__7574 (
            .O(N__37085),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__7573 (
            .O(N__37082),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__7572 (
            .O(N__37079),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__7571 (
            .O(N__37076),
            .I(N__37073));
    LocalMux I__7570 (
            .O(N__37073),
            .I(N__37070));
    Odrv4 I__7569 (
            .O(N__37070),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__7568 (
            .O(N__37067),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__7567 (
            .O(N__37064),
            .I(N__37061));
    LocalMux I__7566 (
            .O(N__37061),
            .I(N__37058));
    Span4Mux_h I__7565 (
            .O(N__37058),
            .I(N__37055));
    Odrv4 I__7564 (
            .O(N__37055),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__7563 (
            .O(N__37052),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    InMux I__7562 (
            .O(N__37049),
            .I(N__37046));
    LocalMux I__7561 (
            .O(N__37046),
            .I(N__37043));
    Odrv4 I__7560 (
            .O(N__37043),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__7559 (
            .O(N__37040),
            .I(bfn_14_16_0_));
    InMux I__7558 (
            .O(N__37037),
            .I(N__37034));
    LocalMux I__7557 (
            .O(N__37034),
            .I(N__37031));
    Odrv4 I__7556 (
            .O(N__37031),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__7555 (
            .O(N__37028),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    InMux I__7554 (
            .O(N__37025),
            .I(N__37022));
    LocalMux I__7553 (
            .O(N__37022),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__7552 (
            .O(N__37019),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__7551 (
            .O(N__37016),
            .I(N__37013));
    LocalMux I__7550 (
            .O(N__37013),
            .I(N__37010));
    Span4Mux_v I__7549 (
            .O(N__37010),
            .I(N__37007));
    Odrv4 I__7548 (
            .O(N__37007),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__7547 (
            .O(N__37004),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    InMux I__7546 (
            .O(N__37001),
            .I(N__36998));
    LocalMux I__7545 (
            .O(N__36998),
            .I(N__36995));
    Span4Mux_h I__7544 (
            .O(N__36995),
            .I(N__36992));
    Odrv4 I__7543 (
            .O(N__36992),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__7542 (
            .O(N__36989),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__7541 (
            .O(N__36986),
            .I(N__36983));
    LocalMux I__7540 (
            .O(N__36983),
            .I(N__36980));
    Odrv4 I__7539 (
            .O(N__36980),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__7538 (
            .O(N__36977),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    InMux I__7537 (
            .O(N__36974),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__7536 (
            .O(N__36971),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    CascadeMux I__7535 (
            .O(N__36968),
            .I(N__36965));
    InMux I__7534 (
            .O(N__36965),
            .I(N__36962));
    LocalMux I__7533 (
            .O(N__36962),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__7532 (
            .O(N__36959),
            .I(N__36956));
    LocalMux I__7531 (
            .O(N__36956),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ));
    InMux I__7530 (
            .O(N__36953),
            .I(N__36950));
    LocalMux I__7529 (
            .O(N__36950),
            .I(N__36947));
    Span4Mux_h I__7528 (
            .O(N__36947),
            .I(N__36944));
    Odrv4 I__7527 (
            .O(N__36944),
            .I(\current_shift_inst.un38_control_input_0_s0_3 ));
    InMux I__7526 (
            .O(N__36941),
            .I(\current_shift_inst.un38_control_input_cry_2_s0 ));
    InMux I__7525 (
            .O(N__36938),
            .I(N__36935));
    LocalMux I__7524 (
            .O(N__36935),
            .I(N__36932));
    Odrv4 I__7523 (
            .O(N__36932),
            .I(\current_shift_inst.un38_control_input_0_s0_4 ));
    InMux I__7522 (
            .O(N__36929),
            .I(\current_shift_inst.un38_control_input_cry_3_s0 ));
    InMux I__7521 (
            .O(N__36926),
            .I(N__36923));
    LocalMux I__7520 (
            .O(N__36923),
            .I(N__36920));
    Span4Mux_h I__7519 (
            .O(N__36920),
            .I(N__36917));
    Odrv4 I__7518 (
            .O(N__36917),
            .I(\current_shift_inst.un38_control_input_0_s0_5 ));
    InMux I__7517 (
            .O(N__36914),
            .I(\current_shift_inst.un38_control_input_cry_4_s0 ));
    InMux I__7516 (
            .O(N__36911),
            .I(N__36908));
    LocalMux I__7515 (
            .O(N__36908),
            .I(N__36905));
    Odrv4 I__7514 (
            .O(N__36905),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__7513 (
            .O(N__36902),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__7512 (
            .O(N__36899),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__7511 (
            .O(N__36896),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__7510 (
            .O(N__36893),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__7509 (
            .O(N__36890),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__7508 (
            .O(N__36887),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__7507 (
            .O(N__36884),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    IoInMux I__7506 (
            .O(N__36881),
            .I(N__36871));
    InMux I__7505 (
            .O(N__36880),
            .I(N__36844));
    InMux I__7504 (
            .O(N__36879),
            .I(N__36844));
    InMux I__7503 (
            .O(N__36878),
            .I(N__36844));
    InMux I__7502 (
            .O(N__36877),
            .I(N__36835));
    InMux I__7501 (
            .O(N__36876),
            .I(N__36835));
    InMux I__7500 (
            .O(N__36875),
            .I(N__36835));
    InMux I__7499 (
            .O(N__36874),
            .I(N__36835));
    LocalMux I__7498 (
            .O(N__36871),
            .I(N__36828));
    InMux I__7497 (
            .O(N__36870),
            .I(N__36819));
    InMux I__7496 (
            .O(N__36869),
            .I(N__36819));
    InMux I__7495 (
            .O(N__36868),
            .I(N__36819));
    InMux I__7494 (
            .O(N__36867),
            .I(N__36819));
    InMux I__7493 (
            .O(N__36866),
            .I(N__36810));
    InMux I__7492 (
            .O(N__36865),
            .I(N__36810));
    InMux I__7491 (
            .O(N__36864),
            .I(N__36810));
    InMux I__7490 (
            .O(N__36863),
            .I(N__36810));
    InMux I__7489 (
            .O(N__36862),
            .I(N__36801));
    InMux I__7488 (
            .O(N__36861),
            .I(N__36801));
    InMux I__7487 (
            .O(N__36860),
            .I(N__36801));
    InMux I__7486 (
            .O(N__36859),
            .I(N__36801));
    InMux I__7485 (
            .O(N__36858),
            .I(N__36792));
    InMux I__7484 (
            .O(N__36857),
            .I(N__36792));
    InMux I__7483 (
            .O(N__36856),
            .I(N__36792));
    InMux I__7482 (
            .O(N__36855),
            .I(N__36792));
    InMux I__7481 (
            .O(N__36854),
            .I(N__36783));
    InMux I__7480 (
            .O(N__36853),
            .I(N__36783));
    InMux I__7479 (
            .O(N__36852),
            .I(N__36783));
    InMux I__7478 (
            .O(N__36851),
            .I(N__36783));
    LocalMux I__7477 (
            .O(N__36844),
            .I(N__36778));
    LocalMux I__7476 (
            .O(N__36835),
            .I(N__36778));
    InMux I__7475 (
            .O(N__36834),
            .I(N__36769));
    InMux I__7474 (
            .O(N__36833),
            .I(N__36769));
    InMux I__7473 (
            .O(N__36832),
            .I(N__36769));
    InMux I__7472 (
            .O(N__36831),
            .I(N__36769));
    IoSpan4Mux I__7471 (
            .O(N__36828),
            .I(N__36766));
    LocalMux I__7470 (
            .O(N__36819),
            .I(N__36761));
    LocalMux I__7469 (
            .O(N__36810),
            .I(N__36761));
    LocalMux I__7468 (
            .O(N__36801),
            .I(N__36750));
    LocalMux I__7467 (
            .O(N__36792),
            .I(N__36750));
    LocalMux I__7466 (
            .O(N__36783),
            .I(N__36750));
    Span4Mux_v I__7465 (
            .O(N__36778),
            .I(N__36750));
    LocalMux I__7464 (
            .O(N__36769),
            .I(N__36750));
    Span4Mux_s2_v I__7463 (
            .O(N__36766),
            .I(N__36747));
    Span4Mux_v I__7462 (
            .O(N__36761),
            .I(N__36742));
    Span4Mux_v I__7461 (
            .O(N__36750),
            .I(N__36742));
    Span4Mux_v I__7460 (
            .O(N__36747),
            .I(N__36739));
    Span4Mux_h I__7459 (
            .O(N__36742),
            .I(N__36736));
    Sp12to4 I__7458 (
            .O(N__36739),
            .I(N__36733));
    Odrv4 I__7457 (
            .O(N__36736),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__7456 (
            .O(N__36733),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__7455 (
            .O(N__36728),
            .I(N__36725));
    LocalMux I__7454 (
            .O(N__36725),
            .I(N__36721));
    InMux I__7453 (
            .O(N__36724),
            .I(N__36718));
    Span4Mux_h I__7452 (
            .O(N__36721),
            .I(N__36715));
    LocalMux I__7451 (
            .O(N__36718),
            .I(N__36712));
    Span4Mux_h I__7450 (
            .O(N__36715),
            .I(N__36709));
    Span12Mux_s10_v I__7449 (
            .O(N__36712),
            .I(N__36706));
    Odrv4 I__7448 (
            .O(N__36709),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    Odrv12 I__7447 (
            .O(N__36706),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__7446 (
            .O(N__36701),
            .I(N__36697));
    InMux I__7445 (
            .O(N__36700),
            .I(N__36693));
    InMux I__7444 (
            .O(N__36697),
            .I(N__36689));
    InMux I__7443 (
            .O(N__36696),
            .I(N__36686));
    LocalMux I__7442 (
            .O(N__36693),
            .I(N__36683));
    InMux I__7441 (
            .O(N__36692),
            .I(N__36679));
    LocalMux I__7440 (
            .O(N__36689),
            .I(N__36676));
    LocalMux I__7439 (
            .O(N__36686),
            .I(N__36673));
    Span4Mux_v I__7438 (
            .O(N__36683),
            .I(N__36670));
    InMux I__7437 (
            .O(N__36682),
            .I(N__36667));
    LocalMux I__7436 (
            .O(N__36679),
            .I(N__36664));
    Span4Mux_h I__7435 (
            .O(N__36676),
            .I(N__36661));
    Span4Mux_h I__7434 (
            .O(N__36673),
            .I(N__36658));
    Span4Mux_h I__7433 (
            .O(N__36670),
            .I(N__36655));
    LocalMux I__7432 (
            .O(N__36667),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__7431 (
            .O(N__36664),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__7430 (
            .O(N__36661),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__7429 (
            .O(N__36658),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__7428 (
            .O(N__36655),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__7427 (
            .O(N__36644),
            .I(bfn_14_12_0_));
    CascadeMux I__7426 (
            .O(N__36641),
            .I(N__36638));
    InMux I__7425 (
            .O(N__36638),
            .I(N__36632));
    InMux I__7424 (
            .O(N__36637),
            .I(N__36632));
    LocalMux I__7423 (
            .O(N__36632),
            .I(N__36628));
    InMux I__7422 (
            .O(N__36631),
            .I(N__36625));
    Span4Mux_h I__7421 (
            .O(N__36628),
            .I(N__36622));
    LocalMux I__7420 (
            .O(N__36625),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__7419 (
            .O(N__36622),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__7418 (
            .O(N__36617),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__7417 (
            .O(N__36614),
            .I(N__36607));
    InMux I__7416 (
            .O(N__36613),
            .I(N__36607));
    InMux I__7415 (
            .O(N__36612),
            .I(N__36604));
    LocalMux I__7414 (
            .O(N__36607),
            .I(N__36601));
    LocalMux I__7413 (
            .O(N__36604),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__7412 (
            .O(N__36601),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__7411 (
            .O(N__36596),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__7410 (
            .O(N__36593),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__7409 (
            .O(N__36590),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__7408 (
            .O(N__36587),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__7407 (
            .O(N__36584),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__7406 (
            .O(N__36581),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__7405 (
            .O(N__36578),
            .I(bfn_14_13_0_));
    InMux I__7404 (
            .O(N__36575),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__7403 (
            .O(N__36572),
            .I(bfn_14_11_0_));
    InMux I__7402 (
            .O(N__36569),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__7401 (
            .O(N__36566),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__7400 (
            .O(N__36563),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__7399 (
            .O(N__36560),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__7398 (
            .O(N__36557),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__7397 (
            .O(N__36554),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__7396 (
            .O(N__36551),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__7395 (
            .O(N__36548),
            .I(N__36545));
    LocalMux I__7394 (
            .O(N__36545),
            .I(N__36542));
    Span4Mux_h I__7393 (
            .O(N__36542),
            .I(N__36539));
    Span4Mux_v I__7392 (
            .O(N__36539),
            .I(N__36536));
    Span4Mux_h I__7391 (
            .O(N__36536),
            .I(N__36533));
    Odrv4 I__7390 (
            .O(N__36533),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    InMux I__7389 (
            .O(N__36530),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__7388 (
            .O(N__36527),
            .I(N__36524));
    InMux I__7387 (
            .O(N__36524),
            .I(N__36521));
    LocalMux I__7386 (
            .O(N__36521),
            .I(N__36518));
    Span4Mux_h I__7385 (
            .O(N__36518),
            .I(N__36515));
    Span4Mux_h I__7384 (
            .O(N__36515),
            .I(N__36512));
    Sp12to4 I__7383 (
            .O(N__36512),
            .I(N__36509));
    Odrv12 I__7382 (
            .O(N__36509),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ));
    InMux I__7381 (
            .O(N__36506),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__7380 (
            .O(N__36503),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__7379 (
            .O(N__36500),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__7378 (
            .O(N__36497),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__7377 (
            .O(N__36494),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    CascadeMux I__7376 (
            .O(N__36491),
            .I(elapsed_time_ns_1_RNI68CN9_0_19_cascade_));
    CascadeMux I__7375 (
            .O(N__36488),
            .I(N__36484));
    InMux I__7374 (
            .O(N__36487),
            .I(N__36481));
    InMux I__7373 (
            .O(N__36484),
            .I(N__36478));
    LocalMux I__7372 (
            .O(N__36481),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    LocalMux I__7371 (
            .O(N__36478),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__7370 (
            .O(N__36473),
            .I(elapsed_time_ns_1_RNI24CN9_0_15_cascade_));
    InMux I__7369 (
            .O(N__36470),
            .I(N__36467));
    LocalMux I__7368 (
            .O(N__36467),
            .I(N__36464));
    Odrv12 I__7367 (
            .O(N__36464),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__7366 (
            .O(N__36461),
            .I(N__36456));
    InMux I__7365 (
            .O(N__36460),
            .I(N__36453));
    InMux I__7364 (
            .O(N__36459),
            .I(N__36450));
    LocalMux I__7363 (
            .O(N__36456),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__7362 (
            .O(N__36453),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__7361 (
            .O(N__36450),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__7360 (
            .O(N__36443),
            .I(N__36437));
    InMux I__7359 (
            .O(N__36442),
            .I(N__36437));
    LocalMux I__7358 (
            .O(N__36437),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__7357 (
            .O(N__36434),
            .I(N__36430));
    InMux I__7356 (
            .O(N__36433),
            .I(N__36427));
    LocalMux I__7355 (
            .O(N__36430),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    LocalMux I__7354 (
            .O(N__36427),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    CascadeMux I__7353 (
            .O(N__36422),
            .I(N__36419));
    InMux I__7352 (
            .O(N__36419),
            .I(N__36413));
    InMux I__7351 (
            .O(N__36418),
            .I(N__36413));
    LocalMux I__7350 (
            .O(N__36413),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__7349 (
            .O(N__36410),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    CascadeMux I__7348 (
            .O(N__36407),
            .I(N__36404));
    InMux I__7347 (
            .O(N__36404),
            .I(N__36401));
    LocalMux I__7346 (
            .O(N__36401),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    InMux I__7345 (
            .O(N__36398),
            .I(N__36392));
    InMux I__7344 (
            .O(N__36397),
            .I(N__36392));
    LocalMux I__7343 (
            .O(N__36392),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    InMux I__7342 (
            .O(N__36389),
            .I(N__36386));
    LocalMux I__7341 (
            .O(N__36386),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    InMux I__7340 (
            .O(N__36383),
            .I(N__36379));
    InMux I__7339 (
            .O(N__36382),
            .I(N__36376));
    LocalMux I__7338 (
            .O(N__36379),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    LocalMux I__7337 (
            .O(N__36376),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    InMux I__7336 (
            .O(N__36371),
            .I(N__36367));
    InMux I__7335 (
            .O(N__36370),
            .I(N__36364));
    LocalMux I__7334 (
            .O(N__36367),
            .I(N__36359));
    LocalMux I__7333 (
            .O(N__36364),
            .I(N__36359));
    Odrv12 I__7332 (
            .O(N__36359),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    InMux I__7331 (
            .O(N__36356),
            .I(N__36353));
    LocalMux I__7330 (
            .O(N__36353),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    InMux I__7329 (
            .O(N__36350),
            .I(N__36347));
    LocalMux I__7328 (
            .O(N__36347),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    CascadeMux I__7327 (
            .O(N__36344),
            .I(N__36340));
    InMux I__7326 (
            .O(N__36343),
            .I(N__36337));
    InMux I__7325 (
            .O(N__36340),
            .I(N__36334));
    LocalMux I__7324 (
            .O(N__36337),
            .I(N__36331));
    LocalMux I__7323 (
            .O(N__36334),
            .I(N__36328));
    Span4Mux_v I__7322 (
            .O(N__36331),
            .I(N__36325));
    Odrv4 I__7321 (
            .O(N__36328),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    Odrv4 I__7320 (
            .O(N__36325),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    InMux I__7319 (
            .O(N__36320),
            .I(N__36317));
    LocalMux I__7318 (
            .O(N__36317),
            .I(N__36313));
    InMux I__7317 (
            .O(N__36316),
            .I(N__36310));
    Odrv4 I__7316 (
            .O(N__36313),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    LocalMux I__7315 (
            .O(N__36310),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__7314 (
            .O(N__36305),
            .I(N__36302));
    InMux I__7313 (
            .O(N__36302),
            .I(N__36299));
    LocalMux I__7312 (
            .O(N__36299),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    InMux I__7311 (
            .O(N__36296),
            .I(N__36293));
    LocalMux I__7310 (
            .O(N__36293),
            .I(N__36289));
    InMux I__7309 (
            .O(N__36292),
            .I(N__36286));
    Odrv4 I__7308 (
            .O(N__36289),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    LocalMux I__7307 (
            .O(N__36286),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__7306 (
            .O(N__36281),
            .I(N__36278));
    InMux I__7305 (
            .O(N__36278),
            .I(N__36275));
    LocalMux I__7304 (
            .O(N__36275),
            .I(N__36272));
    Odrv12 I__7303 (
            .O(N__36272),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    CascadeMux I__7302 (
            .O(N__36269),
            .I(N__36266));
    InMux I__7301 (
            .O(N__36266),
            .I(N__36263));
    LocalMux I__7300 (
            .O(N__36263),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__7299 (
            .O(N__36260),
            .I(N__36257));
    InMux I__7298 (
            .O(N__36257),
            .I(N__36254));
    LocalMux I__7297 (
            .O(N__36254),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    InMux I__7296 (
            .O(N__36251),
            .I(N__36248));
    LocalMux I__7295 (
            .O(N__36248),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    InMux I__7294 (
            .O(N__36245),
            .I(N__36242));
    LocalMux I__7293 (
            .O(N__36242),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__7292 (
            .O(N__36239),
            .I(N__36236));
    LocalMux I__7291 (
            .O(N__36236),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__7290 (
            .O(N__36233),
            .I(N__36230));
    InMux I__7289 (
            .O(N__36230),
            .I(N__36227));
    LocalMux I__7288 (
            .O(N__36227),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__7287 (
            .O(N__36224),
            .I(N__36221));
    InMux I__7286 (
            .O(N__36221),
            .I(N__36218));
    LocalMux I__7285 (
            .O(N__36218),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__7284 (
            .O(N__36215),
            .I(N__36212));
    InMux I__7283 (
            .O(N__36212),
            .I(N__36209));
    LocalMux I__7282 (
            .O(N__36209),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__7281 (
            .O(N__36206),
            .I(N__36203));
    InMux I__7280 (
            .O(N__36203),
            .I(N__36200));
    LocalMux I__7279 (
            .O(N__36200),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__7278 (
            .O(N__36197),
            .I(N__36194));
    InMux I__7277 (
            .O(N__36194),
            .I(N__36191));
    LocalMux I__7276 (
            .O(N__36191),
            .I(N__36188));
    Odrv4 I__7275 (
            .O(N__36188),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__7274 (
            .O(N__36185),
            .I(N__36182));
    InMux I__7273 (
            .O(N__36182),
            .I(N__36179));
    LocalMux I__7272 (
            .O(N__36179),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__7271 (
            .O(N__36176),
            .I(N__36173));
    InMux I__7270 (
            .O(N__36173),
            .I(N__36170));
    LocalMux I__7269 (
            .O(N__36170),
            .I(N__36167));
    Odrv4 I__7268 (
            .O(N__36167),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__7267 (
            .O(N__36164),
            .I(N__36161));
    InMux I__7266 (
            .O(N__36161),
            .I(N__36158));
    LocalMux I__7265 (
            .O(N__36158),
            .I(N__36153));
    InMux I__7264 (
            .O(N__36157),
            .I(N__36150));
    InMux I__7263 (
            .O(N__36156),
            .I(N__36147));
    Span4Mux_v I__7262 (
            .O(N__36153),
            .I(N__36140));
    LocalMux I__7261 (
            .O(N__36150),
            .I(N__36140));
    LocalMux I__7260 (
            .O(N__36147),
            .I(N__36140));
    Span4Mux_v I__7259 (
            .O(N__36140),
            .I(N__36137));
    Span4Mux_v I__7258 (
            .O(N__36137),
            .I(N__36134));
    Span4Mux_v I__7257 (
            .O(N__36134),
            .I(N__36131));
    Odrv4 I__7256 (
            .O(N__36131),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__7255 (
            .O(N__36128),
            .I(N__36125));
    LocalMux I__7254 (
            .O(N__36125),
            .I(N__36121));
    InMux I__7253 (
            .O(N__36124),
            .I(N__36118));
    Span4Mux_v I__7252 (
            .O(N__36121),
            .I(N__36113));
    LocalMux I__7251 (
            .O(N__36118),
            .I(N__36113));
    Span4Mux_v I__7250 (
            .O(N__36113),
            .I(N__36110));
    Span4Mux_v I__7249 (
            .O(N__36110),
            .I(N__36105));
    InMux I__7248 (
            .O(N__36109),
            .I(N__36100));
    InMux I__7247 (
            .O(N__36108),
            .I(N__36100));
    Span4Mux_v I__7246 (
            .O(N__36105),
            .I(N__36097));
    LocalMux I__7245 (
            .O(N__36100),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__7244 (
            .O(N__36097),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    ClkMux I__7243 (
            .O(N__36092),
            .I(N__36089));
    GlobalMux I__7242 (
            .O(N__36089),
            .I(N__36086));
    gio2CtrlBuf I__7241 (
            .O(N__36086),
            .I(delay_hc_input_c_g));
    CascadeMux I__7240 (
            .O(N__36083),
            .I(N__36080));
    InMux I__7239 (
            .O(N__36080),
            .I(N__36077));
    LocalMux I__7238 (
            .O(N__36077),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__7237 (
            .O(N__36074),
            .I(N__36071));
    InMux I__7236 (
            .O(N__36071),
            .I(N__36068));
    LocalMux I__7235 (
            .O(N__36068),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__7234 (
            .O(N__36065),
            .I(N__36062));
    LocalMux I__7233 (
            .O(N__36062),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__7232 (
            .O(N__36059),
            .I(N__36056));
    InMux I__7231 (
            .O(N__36056),
            .I(N__36053));
    LocalMux I__7230 (
            .O(N__36053),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__7229 (
            .O(N__36050),
            .I(N__36047));
    InMux I__7228 (
            .O(N__36047),
            .I(N__36044));
    LocalMux I__7227 (
            .O(N__36044),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__7226 (
            .O(N__36041),
            .I(N__36038));
    LocalMux I__7225 (
            .O(N__36038),
            .I(N__36035));
    Odrv4 I__7224 (
            .O(N__36035),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__7223 (
            .O(N__36032),
            .I(N__36029));
    InMux I__7222 (
            .O(N__36029),
            .I(N__36026));
    LocalMux I__7221 (
            .O(N__36026),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__7220 (
            .O(N__36023),
            .I(N__36020));
    InMux I__7219 (
            .O(N__36020),
            .I(N__36017));
    LocalMux I__7218 (
            .O(N__36017),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    InMux I__7217 (
            .O(N__36014),
            .I(N__36011));
    LocalMux I__7216 (
            .O(N__36011),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__7215 (
            .O(N__36008),
            .I(N__36005));
    LocalMux I__7214 (
            .O(N__36005),
            .I(\current_shift_inst.control_input_axb_25 ));
    InMux I__7213 (
            .O(N__36002),
            .I(N__35999));
    LocalMux I__7212 (
            .O(N__35999),
            .I(\current_shift_inst.control_input_axb_29 ));
    InMux I__7211 (
            .O(N__35996),
            .I(N__35991));
    InMux I__7210 (
            .O(N__35995),
            .I(N__35988));
    InMux I__7209 (
            .O(N__35994),
            .I(N__35985));
    LocalMux I__7208 (
            .O(N__35991),
            .I(N__35982));
    LocalMux I__7207 (
            .O(N__35988),
            .I(N__35977));
    LocalMux I__7206 (
            .O(N__35985),
            .I(N__35977));
    Span4Mux_h I__7205 (
            .O(N__35982),
            .I(N__35974));
    Span4Mux_h I__7204 (
            .O(N__35977),
            .I(N__35971));
    Odrv4 I__7203 (
            .O(N__35974),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__7202 (
            .O(N__35971),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__7201 (
            .O(N__35966),
            .I(N__35962));
    InMux I__7200 (
            .O(N__35965),
            .I(N__35959));
    LocalMux I__7199 (
            .O(N__35962),
            .I(N__35954));
    LocalMux I__7198 (
            .O(N__35959),
            .I(N__35951));
    InMux I__7197 (
            .O(N__35958),
            .I(N__35946));
    InMux I__7196 (
            .O(N__35957),
            .I(N__35946));
    Span4Mux_v I__7195 (
            .O(N__35954),
            .I(N__35943));
    Span4Mux_h I__7194 (
            .O(N__35951),
            .I(N__35940));
    LocalMux I__7193 (
            .O(N__35946),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__7192 (
            .O(N__35943),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__7191 (
            .O(N__35940),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__7190 (
            .O(N__35933),
            .I(N__35930));
    GlobalMux I__7189 (
            .O(N__35930),
            .I(N__35927));
    gio2CtrlBuf I__7188 (
            .O(N__35927),
            .I(delay_tr_input_c_g));
    IoInMux I__7187 (
            .O(N__35924),
            .I(N__35921));
    LocalMux I__7186 (
            .O(N__35921),
            .I(N__35918));
    Span4Mux_s0_v I__7185 (
            .O(N__35918),
            .I(N__35915));
    Span4Mux_v I__7184 (
            .O(N__35915),
            .I(N__35912));
    Span4Mux_v I__7183 (
            .O(N__35912),
            .I(N__35907));
    InMux I__7182 (
            .O(N__35911),
            .I(N__35904));
    InMux I__7181 (
            .O(N__35910),
            .I(N__35901));
    Odrv4 I__7180 (
            .O(N__35907),
            .I(s1_phy_c));
    LocalMux I__7179 (
            .O(N__35904),
            .I(s1_phy_c));
    LocalMux I__7178 (
            .O(N__35901),
            .I(s1_phy_c));
    InMux I__7177 (
            .O(N__35894),
            .I(N__35891));
    LocalMux I__7176 (
            .O(N__35891),
            .I(N__35883));
    InMux I__7175 (
            .O(N__35890),
            .I(N__35878));
    InMux I__7174 (
            .O(N__35889),
            .I(N__35878));
    InMux I__7173 (
            .O(N__35888),
            .I(N__35875));
    CascadeMux I__7172 (
            .O(N__35887),
            .I(N__35871));
    InMux I__7171 (
            .O(N__35886),
            .I(N__35868));
    Span4Mux_v I__7170 (
            .O(N__35883),
            .I(N__35863));
    LocalMux I__7169 (
            .O(N__35878),
            .I(N__35863));
    LocalMux I__7168 (
            .O(N__35875),
            .I(N__35860));
    InMux I__7167 (
            .O(N__35874),
            .I(N__35857));
    InMux I__7166 (
            .O(N__35871),
            .I(N__35854));
    LocalMux I__7165 (
            .O(N__35868),
            .I(N__35851));
    Span4Mux_v I__7164 (
            .O(N__35863),
            .I(N__35848));
    Span4Mux_v I__7163 (
            .O(N__35860),
            .I(N__35845));
    LocalMux I__7162 (
            .O(N__35857),
            .I(state_3));
    LocalMux I__7161 (
            .O(N__35854),
            .I(state_3));
    Odrv12 I__7160 (
            .O(N__35851),
            .I(state_3));
    Odrv4 I__7159 (
            .O(N__35848),
            .I(state_3));
    Odrv4 I__7158 (
            .O(N__35845),
            .I(state_3));
    IoInMux I__7157 (
            .O(N__35834),
            .I(N__35831));
    LocalMux I__7156 (
            .O(N__35831),
            .I(N__35828));
    Odrv12 I__7155 (
            .O(N__35828),
            .I(\current_shift_inst.timer_s1.N_161_i ));
    InMux I__7154 (
            .O(N__35825),
            .I(N__35821));
    InMux I__7153 (
            .O(N__35824),
            .I(N__35818));
    LocalMux I__7152 (
            .O(N__35821),
            .I(N__35815));
    LocalMux I__7151 (
            .O(N__35818),
            .I(N__35811));
    Span4Mux_v I__7150 (
            .O(N__35815),
            .I(N__35808));
    InMux I__7149 (
            .O(N__35814),
            .I(N__35805));
    Span12Mux_s6_v I__7148 (
            .O(N__35811),
            .I(N__35802));
    Span4Mux_v I__7147 (
            .O(N__35808),
            .I(N__35799));
    LocalMux I__7146 (
            .O(N__35805),
            .I(N__35795));
    Span12Mux_v I__7145 (
            .O(N__35802),
            .I(N__35792));
    Span4Mux_v I__7144 (
            .O(N__35799),
            .I(N__35789));
    InMux I__7143 (
            .O(N__35798),
            .I(N__35786));
    Span4Mux_h I__7142 (
            .O(N__35795),
            .I(N__35783));
    Odrv12 I__7141 (
            .O(N__35792),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__7140 (
            .O(N__35789),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__7139 (
            .O(N__35786),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__7138 (
            .O(N__35783),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__7137 (
            .O(N__35774),
            .I(N__35771));
    LocalMux I__7136 (
            .O(N__35771),
            .I(N__35768));
    Odrv4 I__7135 (
            .O(N__35768),
            .I(s2_phy_c));
    InMux I__7134 (
            .O(N__35765),
            .I(N__35762));
    LocalMux I__7133 (
            .O(N__35762),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__7132 (
            .O(N__35759),
            .I(N__35756));
    LocalMux I__7131 (
            .O(N__35756),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__7130 (
            .O(N__35753),
            .I(N__35750));
    LocalMux I__7129 (
            .O(N__35750),
            .I(\current_shift_inst.control_input_axb_18 ));
    InMux I__7128 (
            .O(N__35747),
            .I(N__35744));
    LocalMux I__7127 (
            .O(N__35744),
            .I(\current_shift_inst.control_input_axb_17 ));
    InMux I__7126 (
            .O(N__35741),
            .I(N__35738));
    LocalMux I__7125 (
            .O(N__35738),
            .I(\current_shift_inst.control_input_axb_20 ));
    InMux I__7124 (
            .O(N__35735),
            .I(N__35732));
    LocalMux I__7123 (
            .O(N__35732),
            .I(\current_shift_inst.control_input_axb_21 ));
    InMux I__7122 (
            .O(N__35729),
            .I(N__35726));
    LocalMux I__7121 (
            .O(N__35726),
            .I(\current_shift_inst.control_input_axb_22 ));
    InMux I__7120 (
            .O(N__35723),
            .I(N__35720));
    LocalMux I__7119 (
            .O(N__35720),
            .I(\current_shift_inst.control_input_axb_27 ));
    InMux I__7118 (
            .O(N__35717),
            .I(N__35714));
    LocalMux I__7117 (
            .O(N__35714),
            .I(\current_shift_inst.control_input_axb_26 ));
    InMux I__7116 (
            .O(N__35711),
            .I(N__35708));
    LocalMux I__7115 (
            .O(N__35708),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__7114 (
            .O(N__35705),
            .I(N__35701));
    InMux I__7113 (
            .O(N__35704),
            .I(N__35696));
    LocalMux I__7112 (
            .O(N__35701),
            .I(N__35693));
    InMux I__7111 (
            .O(N__35700),
            .I(N__35690));
    InMux I__7110 (
            .O(N__35699),
            .I(N__35687));
    LocalMux I__7109 (
            .O(N__35696),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__7108 (
            .O(N__35693),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__7107 (
            .O(N__35690),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__7106 (
            .O(N__35687),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__7105 (
            .O(N__35678),
            .I(N__35675));
    LocalMux I__7104 (
            .O(N__35675),
            .I(N__35672));
    Span4Mux_v I__7103 (
            .O(N__35672),
            .I(N__35668));
    InMux I__7102 (
            .O(N__35671),
            .I(N__35664));
    Span4Mux_v I__7101 (
            .O(N__35668),
            .I(N__35660));
    InMux I__7100 (
            .O(N__35667),
            .I(N__35657));
    LocalMux I__7099 (
            .O(N__35664),
            .I(N__35654));
    InMux I__7098 (
            .O(N__35663),
            .I(N__35651));
    Span4Mux_v I__7097 (
            .O(N__35660),
            .I(N__35646));
    LocalMux I__7096 (
            .O(N__35657),
            .I(N__35646));
    Span12Mux_h I__7095 (
            .O(N__35654),
            .I(N__35643));
    LocalMux I__7094 (
            .O(N__35651),
            .I(N__35640));
    Span4Mux_v I__7093 (
            .O(N__35646),
            .I(N__35637));
    Span12Mux_v I__7092 (
            .O(N__35643),
            .I(N__35634));
    Span12Mux_h I__7091 (
            .O(N__35640),
            .I(N__35631));
    Span4Mux_h I__7090 (
            .O(N__35637),
            .I(N__35628));
    Odrv12 I__7089 (
            .O(N__35634),
            .I(il_max_comp1_c));
    Odrv12 I__7088 (
            .O(N__35631),
            .I(il_max_comp1_c));
    Odrv4 I__7087 (
            .O(N__35628),
            .I(il_max_comp1_c));
    IoInMux I__7086 (
            .O(N__35621),
            .I(N__35618));
    LocalMux I__7085 (
            .O(N__35618),
            .I(N__35615));
    Span4Mux_s1_v I__7084 (
            .O(N__35615),
            .I(N__35612));
    Sp12to4 I__7083 (
            .O(N__35612),
            .I(N__35609));
    Span12Mux_h I__7082 (
            .O(N__35609),
            .I(N__35606));
    Span12Mux_v I__7081 (
            .O(N__35606),
            .I(N__35602));
    InMux I__7080 (
            .O(N__35605),
            .I(N__35599));
    Odrv12 I__7079 (
            .O(N__35602),
            .I(test_c));
    LocalMux I__7078 (
            .O(N__35599),
            .I(test_c));
    InMux I__7077 (
            .O(N__35594),
            .I(N__35591));
    LocalMux I__7076 (
            .O(N__35591),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__7075 (
            .O(N__35588),
            .I(N__35585));
    LocalMux I__7074 (
            .O(N__35585),
            .I(\current_shift_inst.control_input_axb_16 ));
    InMux I__7073 (
            .O(N__35582),
            .I(N__35579));
    LocalMux I__7072 (
            .O(N__35579),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__7071 (
            .O(N__35576),
            .I(N__35573));
    LocalMux I__7070 (
            .O(N__35573),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__7069 (
            .O(N__35570),
            .I(N__35567));
    LocalMux I__7068 (
            .O(N__35567),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__7067 (
            .O(N__35564),
            .I(N__35561));
    LocalMux I__7066 (
            .O(N__35561),
            .I(\current_shift_inst.control_input_axb_4 ));
    CascadeMux I__7065 (
            .O(N__35558),
            .I(N__35554));
    CascadeMux I__7064 (
            .O(N__35557),
            .I(N__35551));
    InMux I__7063 (
            .O(N__35554),
            .I(N__35546));
    InMux I__7062 (
            .O(N__35551),
            .I(N__35546));
    LocalMux I__7061 (
            .O(N__35546),
            .I(N__35542));
    InMux I__7060 (
            .O(N__35545),
            .I(N__35539));
    Span4Mux_h I__7059 (
            .O(N__35542),
            .I(N__35536));
    LocalMux I__7058 (
            .O(N__35539),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__7057 (
            .O(N__35536),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__7056 (
            .O(N__35531),
            .I(N__35528));
    LocalMux I__7055 (
            .O(N__35528),
            .I(N__35522));
    InMux I__7054 (
            .O(N__35527),
            .I(N__35519));
    CascadeMux I__7053 (
            .O(N__35526),
            .I(N__35516));
    InMux I__7052 (
            .O(N__35525),
            .I(N__35513));
    Span4Mux_v I__7051 (
            .O(N__35522),
            .I(N__35508));
    LocalMux I__7050 (
            .O(N__35519),
            .I(N__35508));
    InMux I__7049 (
            .O(N__35516),
            .I(N__35505));
    LocalMux I__7048 (
            .O(N__35513),
            .I(N__35502));
    Span4Mux_h I__7047 (
            .O(N__35508),
            .I(N__35499));
    LocalMux I__7046 (
            .O(N__35505),
            .I(N__35496));
    Span4Mux_v I__7045 (
            .O(N__35502),
            .I(N__35493));
    Span4Mux_v I__7044 (
            .O(N__35499),
            .I(N__35488));
    Span4Mux_v I__7043 (
            .O(N__35496),
            .I(N__35488));
    Odrv4 I__7042 (
            .O(N__35493),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__7041 (
            .O(N__35488),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__7040 (
            .O(N__35483),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__7039 (
            .O(N__35480),
            .I(N__35476));
    CascadeMux I__7038 (
            .O(N__35479),
            .I(N__35473));
    InMux I__7037 (
            .O(N__35476),
            .I(N__35470));
    InMux I__7036 (
            .O(N__35473),
            .I(N__35467));
    LocalMux I__7035 (
            .O(N__35470),
            .I(N__35464));
    LocalMux I__7034 (
            .O(N__35467),
            .I(N__35460));
    Span4Mux_h I__7033 (
            .O(N__35464),
            .I(N__35457));
    InMux I__7032 (
            .O(N__35463),
            .I(N__35454));
    Span4Mux_v I__7031 (
            .O(N__35460),
            .I(N__35451));
    Span4Mux_h I__7030 (
            .O(N__35457),
            .I(N__35448));
    LocalMux I__7029 (
            .O(N__35454),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__7028 (
            .O(N__35451),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__7027 (
            .O(N__35448),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__7026 (
            .O(N__35441),
            .I(N__35437));
    InMux I__7025 (
            .O(N__35440),
            .I(N__35434));
    LocalMux I__7024 (
            .O(N__35437),
            .I(N__35431));
    LocalMux I__7023 (
            .O(N__35434),
            .I(N__35426));
    Span4Mux_v I__7022 (
            .O(N__35431),
            .I(N__35423));
    InMux I__7021 (
            .O(N__35430),
            .I(N__35418));
    InMux I__7020 (
            .O(N__35429),
            .I(N__35418));
    Span4Mux_v I__7019 (
            .O(N__35426),
            .I(N__35415));
    Sp12to4 I__7018 (
            .O(N__35423),
            .I(N__35410));
    LocalMux I__7017 (
            .O(N__35418),
            .I(N__35410));
    Span4Mux_v I__7016 (
            .O(N__35415),
            .I(N__35407));
    Odrv12 I__7015 (
            .O(N__35410),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__7014 (
            .O(N__35407),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__7013 (
            .O(N__35402),
            .I(bfn_13_13_0_));
    InMux I__7012 (
            .O(N__35399),
            .I(N__35395));
    InMux I__7011 (
            .O(N__35398),
            .I(N__35392));
    LocalMux I__7010 (
            .O(N__35395),
            .I(N__35386));
    LocalMux I__7009 (
            .O(N__35392),
            .I(N__35386));
    InMux I__7008 (
            .O(N__35391),
            .I(N__35383));
    Span4Mux_v I__7007 (
            .O(N__35386),
            .I(N__35380));
    LocalMux I__7006 (
            .O(N__35383),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__7005 (
            .O(N__35380),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__7004 (
            .O(N__35375),
            .I(N__35371));
    InMux I__7003 (
            .O(N__35374),
            .I(N__35367));
    LocalMux I__7002 (
            .O(N__35371),
            .I(N__35364));
    InMux I__7001 (
            .O(N__35370),
            .I(N__35360));
    LocalMux I__7000 (
            .O(N__35367),
            .I(N__35357));
    Span4Mux_v I__6999 (
            .O(N__35364),
            .I(N__35354));
    InMux I__6998 (
            .O(N__35363),
            .I(N__35351));
    LocalMux I__6997 (
            .O(N__35360),
            .I(N__35348));
    Span4Mux_v I__6996 (
            .O(N__35357),
            .I(N__35345));
    Span4Mux_v I__6995 (
            .O(N__35354),
            .I(N__35342));
    LocalMux I__6994 (
            .O(N__35351),
            .I(N__35337));
    Span12Mux_v I__6993 (
            .O(N__35348),
            .I(N__35337));
    Span4Mux_h I__6992 (
            .O(N__35345),
            .I(N__35334));
    Span4Mux_h I__6991 (
            .O(N__35342),
            .I(N__35331));
    Odrv12 I__6990 (
            .O(N__35337),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__6989 (
            .O(N__35334),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__6988 (
            .O(N__35331),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__6987 (
            .O(N__35324),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__6986 (
            .O(N__35321),
            .I(N__35318));
    LocalMux I__6985 (
            .O(N__35318),
            .I(N__35314));
    InMux I__6984 (
            .O(N__35317),
            .I(N__35311));
    Span4Mux_h I__6983 (
            .O(N__35314),
            .I(N__35308));
    LocalMux I__6982 (
            .O(N__35311),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv4 I__6981 (
            .O(N__35308),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__6980 (
            .O(N__35303),
            .I(N__35300));
    InMux I__6979 (
            .O(N__35300),
            .I(N__35296));
    InMux I__6978 (
            .O(N__35299),
            .I(N__35293));
    LocalMux I__6977 (
            .O(N__35296),
            .I(N__35287));
    LocalMux I__6976 (
            .O(N__35293),
            .I(N__35287));
    InMux I__6975 (
            .O(N__35292),
            .I(N__35284));
    Span4Mux_h I__6974 (
            .O(N__35287),
            .I(N__35281));
    LocalMux I__6973 (
            .O(N__35284),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__6972 (
            .O(N__35281),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__6971 (
            .O(N__35276),
            .I(N__35272));
    InMux I__6970 (
            .O(N__35275),
            .I(N__35267));
    LocalMux I__6969 (
            .O(N__35272),
            .I(N__35264));
    InMux I__6968 (
            .O(N__35271),
            .I(N__35259));
    InMux I__6967 (
            .O(N__35270),
            .I(N__35259));
    LocalMux I__6966 (
            .O(N__35267),
            .I(N__35256));
    Span4Mux_v I__6965 (
            .O(N__35264),
            .I(N__35251));
    LocalMux I__6964 (
            .O(N__35259),
            .I(N__35251));
    Span4Mux_h I__6963 (
            .O(N__35256),
            .I(N__35248));
    Span4Mux_h I__6962 (
            .O(N__35251),
            .I(N__35243));
    Span4Mux_v I__6961 (
            .O(N__35248),
            .I(N__35243));
    Odrv4 I__6960 (
            .O(N__35243),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__6959 (
            .O(N__35240),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__6958 (
            .O(N__35237),
            .I(N__35234));
    LocalMux I__6957 (
            .O(N__35234),
            .I(N__35230));
    InMux I__6956 (
            .O(N__35233),
            .I(N__35227));
    Span4Mux_h I__6955 (
            .O(N__35230),
            .I(N__35224));
    LocalMux I__6954 (
            .O(N__35227),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__6953 (
            .O(N__35224),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__6952 (
            .O(N__35219),
            .I(N__35215));
    CascadeMux I__6951 (
            .O(N__35218),
            .I(N__35212));
    InMux I__6950 (
            .O(N__35215),
            .I(N__35207));
    InMux I__6949 (
            .O(N__35212),
            .I(N__35207));
    LocalMux I__6948 (
            .O(N__35207),
            .I(N__35203));
    InMux I__6947 (
            .O(N__35206),
            .I(N__35200));
    Span4Mux_h I__6946 (
            .O(N__35203),
            .I(N__35197));
    LocalMux I__6945 (
            .O(N__35200),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__6944 (
            .O(N__35197),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__6943 (
            .O(N__35192),
            .I(N__35186));
    InMux I__6942 (
            .O(N__35191),
            .I(N__35183));
    InMux I__6941 (
            .O(N__35190),
            .I(N__35180));
    InMux I__6940 (
            .O(N__35189),
            .I(N__35177));
    LocalMux I__6939 (
            .O(N__35186),
            .I(N__35170));
    LocalMux I__6938 (
            .O(N__35183),
            .I(N__35170));
    LocalMux I__6937 (
            .O(N__35180),
            .I(N__35170));
    LocalMux I__6936 (
            .O(N__35177),
            .I(N__35167));
    Span4Mux_v I__6935 (
            .O(N__35170),
            .I(N__35164));
    Span4Mux_h I__6934 (
            .O(N__35167),
            .I(N__35161));
    Odrv4 I__6933 (
            .O(N__35164),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__6932 (
            .O(N__35161),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__6931 (
            .O(N__35156),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__6930 (
            .O(N__35153),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__6929 (
            .O(N__35150),
            .I(N__35144));
    InMux I__6928 (
            .O(N__35149),
            .I(N__35141));
    InMux I__6927 (
            .O(N__35148),
            .I(N__35138));
    InMux I__6926 (
            .O(N__35147),
            .I(N__35135));
    LocalMux I__6925 (
            .O(N__35144),
            .I(N__35132));
    LocalMux I__6924 (
            .O(N__35141),
            .I(N__35127));
    LocalMux I__6923 (
            .O(N__35138),
            .I(N__35127));
    LocalMux I__6922 (
            .O(N__35135),
            .I(N__35124));
    Span4Mux_h I__6921 (
            .O(N__35132),
            .I(N__35121));
    Span4Mux_v I__6920 (
            .O(N__35127),
            .I(N__35118));
    Span4Mux_h I__6919 (
            .O(N__35124),
            .I(N__35115));
    Span4Mux_v I__6918 (
            .O(N__35121),
            .I(N__35112));
    Odrv4 I__6917 (
            .O(N__35118),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__6916 (
            .O(N__35115),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__6915 (
            .O(N__35112),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    CEMux I__6914 (
            .O(N__35105),
            .I(N__35101));
    CEMux I__6913 (
            .O(N__35104),
            .I(N__35096));
    LocalMux I__6912 (
            .O(N__35101),
            .I(N__35093));
    CEMux I__6911 (
            .O(N__35100),
            .I(N__35090));
    CEMux I__6910 (
            .O(N__35099),
            .I(N__35087));
    LocalMux I__6909 (
            .O(N__35096),
            .I(N__35083));
    Span4Mux_v I__6908 (
            .O(N__35093),
            .I(N__35080));
    LocalMux I__6907 (
            .O(N__35090),
            .I(N__35077));
    LocalMux I__6906 (
            .O(N__35087),
            .I(N__35074));
    CEMux I__6905 (
            .O(N__35086),
            .I(N__35071));
    Span4Mux_h I__6904 (
            .O(N__35083),
            .I(N__35068));
    Span4Mux_h I__6903 (
            .O(N__35080),
            .I(N__35065));
    Span4Mux_h I__6902 (
            .O(N__35077),
            .I(N__35062));
    Span4Mux_v I__6901 (
            .O(N__35074),
            .I(N__35059));
    LocalMux I__6900 (
            .O(N__35071),
            .I(N__35056));
    Span4Mux_v I__6899 (
            .O(N__35068),
            .I(N__35053));
    Span4Mux_v I__6898 (
            .O(N__35065),
            .I(N__35048));
    Span4Mux_v I__6897 (
            .O(N__35062),
            .I(N__35048));
    Span4Mux_v I__6896 (
            .O(N__35059),
            .I(N__35043));
    Span4Mux_h I__6895 (
            .O(N__35056),
            .I(N__35043));
    Odrv4 I__6894 (
            .O(N__35053),
            .I(\delay_measurement_inst.delay_tr_timer.N_165_i ));
    Odrv4 I__6893 (
            .O(N__35048),
            .I(\delay_measurement_inst.delay_tr_timer.N_165_i ));
    Odrv4 I__6892 (
            .O(N__35043),
            .I(\delay_measurement_inst.delay_tr_timer.N_165_i ));
    InMux I__6891 (
            .O(N__35036),
            .I(N__35030));
    InMux I__6890 (
            .O(N__35035),
            .I(N__35030));
    LocalMux I__6889 (
            .O(N__35030),
            .I(N__35026));
    InMux I__6888 (
            .O(N__35029),
            .I(N__35023));
    Span4Mux_h I__6887 (
            .O(N__35026),
            .I(N__35020));
    LocalMux I__6886 (
            .O(N__35023),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__6885 (
            .O(N__35020),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__6884 (
            .O(N__35015),
            .I(N__35011));
    InMux I__6883 (
            .O(N__35014),
            .I(N__35008));
    LocalMux I__6882 (
            .O(N__35011),
            .I(N__35002));
    LocalMux I__6881 (
            .O(N__35008),
            .I(N__35002));
    InMux I__6880 (
            .O(N__35007),
            .I(N__34999));
    Span4Mux_v I__6879 (
            .O(N__35002),
            .I(N__34993));
    LocalMux I__6878 (
            .O(N__34999),
            .I(N__34993));
    InMux I__6877 (
            .O(N__34998),
            .I(N__34990));
    Span4Mux_h I__6876 (
            .O(N__34993),
            .I(N__34985));
    LocalMux I__6875 (
            .O(N__34990),
            .I(N__34985));
    Odrv4 I__6874 (
            .O(N__34985),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__6873 (
            .O(N__34982),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__6872 (
            .O(N__34979),
            .I(N__34976));
    InMux I__6871 (
            .O(N__34976),
            .I(N__34973));
    LocalMux I__6870 (
            .O(N__34973),
            .I(N__34969));
    InMux I__6869 (
            .O(N__34972),
            .I(N__34966));
    Span4Mux_v I__6868 (
            .O(N__34969),
            .I(N__34962));
    LocalMux I__6867 (
            .O(N__34966),
            .I(N__34959));
    InMux I__6866 (
            .O(N__34965),
            .I(N__34956));
    Span4Mux_h I__6865 (
            .O(N__34962),
            .I(N__34953));
    Span4Mux_h I__6864 (
            .O(N__34959),
            .I(N__34950));
    LocalMux I__6863 (
            .O(N__34956),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__6862 (
            .O(N__34953),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__6861 (
            .O(N__34950),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__6860 (
            .O(N__34943),
            .I(N__34939));
    InMux I__6859 (
            .O(N__34942),
            .I(N__34936));
    LocalMux I__6858 (
            .O(N__34939),
            .I(N__34931));
    LocalMux I__6857 (
            .O(N__34936),
            .I(N__34928));
    InMux I__6856 (
            .O(N__34935),
            .I(N__34925));
    CascadeMux I__6855 (
            .O(N__34934),
            .I(N__34922));
    Span4Mux_h I__6854 (
            .O(N__34931),
            .I(N__34919));
    Span4Mux_v I__6853 (
            .O(N__34928),
            .I(N__34916));
    LocalMux I__6852 (
            .O(N__34925),
            .I(N__34913));
    InMux I__6851 (
            .O(N__34922),
            .I(N__34910));
    Span4Mux_v I__6850 (
            .O(N__34919),
            .I(N__34907));
    Span4Mux_h I__6849 (
            .O(N__34916),
            .I(N__34900));
    Span4Mux_v I__6848 (
            .O(N__34913),
            .I(N__34900));
    LocalMux I__6847 (
            .O(N__34910),
            .I(N__34900));
    Odrv4 I__6846 (
            .O(N__34907),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__6845 (
            .O(N__34900),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__6844 (
            .O(N__34895),
            .I(bfn_13_12_0_));
    CascadeMux I__6843 (
            .O(N__34892),
            .I(N__34888));
    CascadeMux I__6842 (
            .O(N__34891),
            .I(N__34885));
    InMux I__6841 (
            .O(N__34888),
            .I(N__34882));
    InMux I__6840 (
            .O(N__34885),
            .I(N__34879));
    LocalMux I__6839 (
            .O(N__34882),
            .I(N__34875));
    LocalMux I__6838 (
            .O(N__34879),
            .I(N__34872));
    InMux I__6837 (
            .O(N__34878),
            .I(N__34869));
    Span4Mux_v I__6836 (
            .O(N__34875),
            .I(N__34866));
    Span4Mux_h I__6835 (
            .O(N__34872),
            .I(N__34863));
    LocalMux I__6834 (
            .O(N__34869),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__6833 (
            .O(N__34866),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__6832 (
            .O(N__34863),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__6831 (
            .O(N__34856),
            .I(N__34853));
    LocalMux I__6830 (
            .O(N__34853),
            .I(N__34849));
    InMux I__6829 (
            .O(N__34852),
            .I(N__34846));
    Span4Mux_v I__6828 (
            .O(N__34849),
            .I(N__34840));
    LocalMux I__6827 (
            .O(N__34846),
            .I(N__34840));
    InMux I__6826 (
            .O(N__34845),
            .I(N__34837));
    Span4Mux_v I__6825 (
            .O(N__34840),
            .I(N__34834));
    LocalMux I__6824 (
            .O(N__34837),
            .I(N__34831));
    Span4Mux_h I__6823 (
            .O(N__34834),
            .I(N__34825));
    Span4Mux_h I__6822 (
            .O(N__34831),
            .I(N__34825));
    InMux I__6821 (
            .O(N__34830),
            .I(N__34822));
    Span4Mux_v I__6820 (
            .O(N__34825),
            .I(N__34817));
    LocalMux I__6819 (
            .O(N__34822),
            .I(N__34817));
    Odrv4 I__6818 (
            .O(N__34817),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__6817 (
            .O(N__34814),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__6816 (
            .O(N__34811),
            .I(N__34808));
    InMux I__6815 (
            .O(N__34808),
            .I(N__34804));
    InMux I__6814 (
            .O(N__34807),
            .I(N__34801));
    LocalMux I__6813 (
            .O(N__34804),
            .I(N__34795));
    LocalMux I__6812 (
            .O(N__34801),
            .I(N__34795));
    InMux I__6811 (
            .O(N__34800),
            .I(N__34792));
    Span4Mux_h I__6810 (
            .O(N__34795),
            .I(N__34789));
    LocalMux I__6809 (
            .O(N__34792),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__6808 (
            .O(N__34789),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__6807 (
            .O(N__34784),
            .I(N__34781));
    LocalMux I__6806 (
            .O(N__34781),
            .I(N__34778));
    Span4Mux_v I__6805 (
            .O(N__34778),
            .I(N__34773));
    InMux I__6804 (
            .O(N__34777),
            .I(N__34770));
    InMux I__6803 (
            .O(N__34776),
            .I(N__34767));
    Span4Mux_v I__6802 (
            .O(N__34773),
            .I(N__34759));
    LocalMux I__6801 (
            .O(N__34770),
            .I(N__34759));
    LocalMux I__6800 (
            .O(N__34767),
            .I(N__34759));
    InMux I__6799 (
            .O(N__34766),
            .I(N__34756));
    Span4Mux_h I__6798 (
            .O(N__34759),
            .I(N__34751));
    LocalMux I__6797 (
            .O(N__34756),
            .I(N__34751));
    Odrv4 I__6796 (
            .O(N__34751),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__6795 (
            .O(N__34748),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__6794 (
            .O(N__34745),
            .I(N__34742));
    InMux I__6793 (
            .O(N__34742),
            .I(N__34738));
    InMux I__6792 (
            .O(N__34741),
            .I(N__34735));
    LocalMux I__6791 (
            .O(N__34738),
            .I(N__34729));
    LocalMux I__6790 (
            .O(N__34735),
            .I(N__34729));
    InMux I__6789 (
            .O(N__34734),
            .I(N__34726));
    Span4Mux_h I__6788 (
            .O(N__34729),
            .I(N__34723));
    LocalMux I__6787 (
            .O(N__34726),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__6786 (
            .O(N__34723),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__6785 (
            .O(N__34718),
            .I(N__34713));
    InMux I__6784 (
            .O(N__34717),
            .I(N__34710));
    InMux I__6783 (
            .O(N__34716),
            .I(N__34707));
    LocalMux I__6782 (
            .O(N__34713),
            .I(N__34703));
    LocalMux I__6781 (
            .O(N__34710),
            .I(N__34698));
    LocalMux I__6780 (
            .O(N__34707),
            .I(N__34698));
    InMux I__6779 (
            .O(N__34706),
            .I(N__34695));
    Span4Mux_v I__6778 (
            .O(N__34703),
            .I(N__34690));
    Span4Mux_v I__6777 (
            .O(N__34698),
            .I(N__34690));
    LocalMux I__6776 (
            .O(N__34695),
            .I(N__34687));
    Span4Mux_h I__6775 (
            .O(N__34690),
            .I(N__34684));
    Span4Mux_v I__6774 (
            .O(N__34687),
            .I(N__34681));
    Odrv4 I__6773 (
            .O(N__34684),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv4 I__6772 (
            .O(N__34681),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__6771 (
            .O(N__34676),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__6770 (
            .O(N__34673),
            .I(N__34670));
    InMux I__6769 (
            .O(N__34670),
            .I(N__34666));
    InMux I__6768 (
            .O(N__34669),
            .I(N__34663));
    LocalMux I__6767 (
            .O(N__34666),
            .I(N__34657));
    LocalMux I__6766 (
            .O(N__34663),
            .I(N__34657));
    InMux I__6765 (
            .O(N__34662),
            .I(N__34654));
    Span4Mux_h I__6764 (
            .O(N__34657),
            .I(N__34651));
    LocalMux I__6763 (
            .O(N__34654),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__6762 (
            .O(N__34651),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__6761 (
            .O(N__34646),
            .I(N__34641));
    InMux I__6760 (
            .O(N__34645),
            .I(N__34637));
    CascadeMux I__6759 (
            .O(N__34644),
            .I(N__34634));
    LocalMux I__6758 (
            .O(N__34641),
            .I(N__34631));
    InMux I__6757 (
            .O(N__34640),
            .I(N__34628));
    LocalMux I__6756 (
            .O(N__34637),
            .I(N__34625));
    InMux I__6755 (
            .O(N__34634),
            .I(N__34622));
    Span4Mux_h I__6754 (
            .O(N__34631),
            .I(N__34617));
    LocalMux I__6753 (
            .O(N__34628),
            .I(N__34617));
    Span4Mux_h I__6752 (
            .O(N__34625),
            .I(N__34612));
    LocalMux I__6751 (
            .O(N__34622),
            .I(N__34612));
    Span4Mux_h I__6750 (
            .O(N__34617),
            .I(N__34609));
    Span4Mux_v I__6749 (
            .O(N__34612),
            .I(N__34606));
    Odrv4 I__6748 (
            .O(N__34609),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv4 I__6747 (
            .O(N__34606),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__6746 (
            .O(N__34601),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__6745 (
            .O(N__34598),
            .I(N__34592));
    InMux I__6744 (
            .O(N__34597),
            .I(N__34592));
    LocalMux I__6743 (
            .O(N__34592),
            .I(N__34588));
    InMux I__6742 (
            .O(N__34591),
            .I(N__34585));
    Span4Mux_h I__6741 (
            .O(N__34588),
            .I(N__34582));
    LocalMux I__6740 (
            .O(N__34585),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv4 I__6739 (
            .O(N__34582),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__6738 (
            .O(N__34577),
            .I(N__34573));
    InMux I__6737 (
            .O(N__34576),
            .I(N__34570));
    LocalMux I__6736 (
            .O(N__34573),
            .I(N__34567));
    LocalMux I__6735 (
            .O(N__34570),
            .I(N__34562));
    Span4Mux_v I__6734 (
            .O(N__34567),
            .I(N__34559));
    InMux I__6733 (
            .O(N__34566),
            .I(N__34556));
    InMux I__6732 (
            .O(N__34565),
            .I(N__34553));
    Span4Mux_h I__6731 (
            .O(N__34562),
            .I(N__34546));
    Span4Mux_h I__6730 (
            .O(N__34559),
            .I(N__34546));
    LocalMux I__6729 (
            .O(N__34556),
            .I(N__34546));
    LocalMux I__6728 (
            .O(N__34553),
            .I(N__34543));
    Odrv4 I__6727 (
            .O(N__34546),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__6726 (
            .O(N__34543),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__6725 (
            .O(N__34538),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__6724 (
            .O(N__34535),
            .I(N__34529));
    InMux I__6723 (
            .O(N__34534),
            .I(N__34529));
    LocalMux I__6722 (
            .O(N__34529),
            .I(N__34525));
    InMux I__6721 (
            .O(N__34528),
            .I(N__34522));
    Span4Mux_h I__6720 (
            .O(N__34525),
            .I(N__34519));
    LocalMux I__6719 (
            .O(N__34522),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__6718 (
            .O(N__34519),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__6717 (
            .O(N__34514),
            .I(N__34509));
    InMux I__6716 (
            .O(N__34513),
            .I(N__34505));
    InMux I__6715 (
            .O(N__34512),
            .I(N__34502));
    LocalMux I__6714 (
            .O(N__34509),
            .I(N__34499));
    InMux I__6713 (
            .O(N__34508),
            .I(N__34496));
    LocalMux I__6712 (
            .O(N__34505),
            .I(N__34493));
    LocalMux I__6711 (
            .O(N__34502),
            .I(N__34490));
    Span4Mux_v I__6710 (
            .O(N__34499),
            .I(N__34485));
    LocalMux I__6709 (
            .O(N__34496),
            .I(N__34485));
    Span4Mux_h I__6708 (
            .O(N__34493),
            .I(N__34482));
    Span4Mux_h I__6707 (
            .O(N__34490),
            .I(N__34479));
    Odrv4 I__6706 (
            .O(N__34485),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__6705 (
            .O(N__34482),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__6704 (
            .O(N__34479),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__6703 (
            .O(N__34472),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__6702 (
            .O(N__34469),
            .I(N__34464));
    InMux I__6701 (
            .O(N__34468),
            .I(N__34459));
    InMux I__6700 (
            .O(N__34467),
            .I(N__34459));
    LocalMux I__6699 (
            .O(N__34464),
            .I(N__34453));
    LocalMux I__6698 (
            .O(N__34459),
            .I(N__34453));
    InMux I__6697 (
            .O(N__34458),
            .I(N__34450));
    Span4Mux_v I__6696 (
            .O(N__34453),
            .I(N__34445));
    LocalMux I__6695 (
            .O(N__34450),
            .I(N__34445));
    Span4Mux_h I__6694 (
            .O(N__34445),
            .I(N__34442));
    Odrv4 I__6693 (
            .O(N__34442),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__6692 (
            .O(N__34439),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__6691 (
            .O(N__34436),
            .I(N__34433));
    InMux I__6690 (
            .O(N__34433),
            .I(N__34430));
    LocalMux I__6689 (
            .O(N__34430),
            .I(N__34425));
    InMux I__6688 (
            .O(N__34429),
            .I(N__34422));
    InMux I__6687 (
            .O(N__34428),
            .I(N__34419));
    Span4Mux_v I__6686 (
            .O(N__34425),
            .I(N__34416));
    LocalMux I__6685 (
            .O(N__34422),
            .I(N__34413));
    LocalMux I__6684 (
            .O(N__34419),
            .I(N__34408));
    Span4Mux_h I__6683 (
            .O(N__34416),
            .I(N__34408));
    Span4Mux_h I__6682 (
            .O(N__34413),
            .I(N__34405));
    Odrv4 I__6681 (
            .O(N__34408),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__6680 (
            .O(N__34405),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    CascadeMux I__6679 (
            .O(N__34400),
            .I(N__34397));
    InMux I__6678 (
            .O(N__34397),
            .I(N__34392));
    InMux I__6677 (
            .O(N__34396),
            .I(N__34389));
    InMux I__6676 (
            .O(N__34395),
            .I(N__34386));
    LocalMux I__6675 (
            .O(N__34392),
            .I(N__34380));
    LocalMux I__6674 (
            .O(N__34389),
            .I(N__34380));
    LocalMux I__6673 (
            .O(N__34386),
            .I(N__34377));
    InMux I__6672 (
            .O(N__34385),
            .I(N__34374));
    Span4Mux_v I__6671 (
            .O(N__34380),
            .I(N__34371));
    Span4Mux_h I__6670 (
            .O(N__34377),
            .I(N__34366));
    LocalMux I__6669 (
            .O(N__34374),
            .I(N__34366));
    Span4Mux_h I__6668 (
            .O(N__34371),
            .I(N__34363));
    Span4Mux_v I__6667 (
            .O(N__34366),
            .I(N__34360));
    Odrv4 I__6666 (
            .O(N__34363),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    Odrv4 I__6665 (
            .O(N__34360),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__6664 (
            .O(N__34355),
            .I(bfn_13_11_0_));
    CascadeMux I__6663 (
            .O(N__34352),
            .I(N__34349));
    InMux I__6662 (
            .O(N__34349),
            .I(N__34344));
    InMux I__6661 (
            .O(N__34348),
            .I(N__34341));
    InMux I__6660 (
            .O(N__34347),
            .I(N__34338));
    LocalMux I__6659 (
            .O(N__34344),
            .I(N__34335));
    LocalMux I__6658 (
            .O(N__34341),
            .I(N__34332));
    LocalMux I__6657 (
            .O(N__34338),
            .I(N__34327));
    Span4Mux_v I__6656 (
            .O(N__34335),
            .I(N__34327));
    Span4Mux_h I__6655 (
            .O(N__34332),
            .I(N__34324));
    Odrv4 I__6654 (
            .O(N__34327),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__6653 (
            .O(N__34324),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    CascadeMux I__6652 (
            .O(N__34319),
            .I(N__34316));
    InMux I__6651 (
            .O(N__34316),
            .I(N__34311));
    InMux I__6650 (
            .O(N__34315),
            .I(N__34308));
    CascadeMux I__6649 (
            .O(N__34314),
            .I(N__34305));
    LocalMux I__6648 (
            .O(N__34311),
            .I(N__34301));
    LocalMux I__6647 (
            .O(N__34308),
            .I(N__34298));
    InMux I__6646 (
            .O(N__34305),
            .I(N__34295));
    InMux I__6645 (
            .O(N__34304),
            .I(N__34292));
    Span4Mux_v I__6644 (
            .O(N__34301),
            .I(N__34285));
    Span4Mux_h I__6643 (
            .O(N__34298),
            .I(N__34285));
    LocalMux I__6642 (
            .O(N__34295),
            .I(N__34285));
    LocalMux I__6641 (
            .O(N__34292),
            .I(N__34282));
    Span4Mux_h I__6640 (
            .O(N__34285),
            .I(N__34279));
    Odrv12 I__6639 (
            .O(N__34282),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__6638 (
            .O(N__34279),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__6637 (
            .O(N__34274),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__6636 (
            .O(N__34271),
            .I(N__34268));
    InMux I__6635 (
            .O(N__34268),
            .I(N__34264));
    InMux I__6634 (
            .O(N__34267),
            .I(N__34261));
    LocalMux I__6633 (
            .O(N__34264),
            .I(N__34255));
    LocalMux I__6632 (
            .O(N__34261),
            .I(N__34255));
    InMux I__6631 (
            .O(N__34260),
            .I(N__34252));
    Span4Mux_h I__6630 (
            .O(N__34255),
            .I(N__34249));
    LocalMux I__6629 (
            .O(N__34252),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__6628 (
            .O(N__34249),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__6627 (
            .O(N__34244),
            .I(N__34240));
    InMux I__6626 (
            .O(N__34243),
            .I(N__34236));
    LocalMux I__6625 (
            .O(N__34240),
            .I(N__34233));
    InMux I__6624 (
            .O(N__34239),
            .I(N__34230));
    LocalMux I__6623 (
            .O(N__34236),
            .I(N__34226));
    Span4Mux_v I__6622 (
            .O(N__34233),
            .I(N__34221));
    LocalMux I__6621 (
            .O(N__34230),
            .I(N__34221));
    InMux I__6620 (
            .O(N__34229),
            .I(N__34218));
    Span4Mux_v I__6619 (
            .O(N__34226),
            .I(N__34215));
    Span4Mux_h I__6618 (
            .O(N__34221),
            .I(N__34210));
    LocalMux I__6617 (
            .O(N__34218),
            .I(N__34210));
    Odrv4 I__6616 (
            .O(N__34215),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__6615 (
            .O(N__34210),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__6614 (
            .O(N__34205),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__6613 (
            .O(N__34202),
            .I(N__34199));
    InMux I__6612 (
            .O(N__34199),
            .I(N__34195));
    InMux I__6611 (
            .O(N__34198),
            .I(N__34192));
    LocalMux I__6610 (
            .O(N__34195),
            .I(N__34186));
    LocalMux I__6609 (
            .O(N__34192),
            .I(N__34186));
    InMux I__6608 (
            .O(N__34191),
            .I(N__34183));
    Span4Mux_h I__6607 (
            .O(N__34186),
            .I(N__34180));
    LocalMux I__6606 (
            .O(N__34183),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__6605 (
            .O(N__34180),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__6604 (
            .O(N__34175),
            .I(N__34170));
    InMux I__6603 (
            .O(N__34174),
            .I(N__34167));
    CascadeMux I__6602 (
            .O(N__34173),
            .I(N__34163));
    LocalMux I__6601 (
            .O(N__34170),
            .I(N__34160));
    LocalMux I__6600 (
            .O(N__34167),
            .I(N__34157));
    InMux I__6599 (
            .O(N__34166),
            .I(N__34154));
    InMux I__6598 (
            .O(N__34163),
            .I(N__34151));
    Span4Mux_h I__6597 (
            .O(N__34160),
            .I(N__34144));
    Span4Mux_h I__6596 (
            .O(N__34157),
            .I(N__34144));
    LocalMux I__6595 (
            .O(N__34154),
            .I(N__34144));
    LocalMux I__6594 (
            .O(N__34151),
            .I(N__34141));
    Odrv4 I__6593 (
            .O(N__34144),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    Odrv4 I__6592 (
            .O(N__34141),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__6591 (
            .O(N__34136),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__6590 (
            .O(N__34133),
            .I(N__34130));
    InMux I__6589 (
            .O(N__34130),
            .I(N__34126));
    InMux I__6588 (
            .O(N__34129),
            .I(N__34123));
    LocalMux I__6587 (
            .O(N__34126),
            .I(N__34117));
    LocalMux I__6586 (
            .O(N__34123),
            .I(N__34117));
    InMux I__6585 (
            .O(N__34122),
            .I(N__34114));
    Span4Mux_h I__6584 (
            .O(N__34117),
            .I(N__34111));
    LocalMux I__6583 (
            .O(N__34114),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__6582 (
            .O(N__34111),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__6581 (
            .O(N__34106),
            .I(N__34103));
    LocalMux I__6580 (
            .O(N__34103),
            .I(N__34097));
    InMux I__6579 (
            .O(N__34102),
            .I(N__34092));
    InMux I__6578 (
            .O(N__34101),
            .I(N__34092));
    InMux I__6577 (
            .O(N__34100),
            .I(N__34089));
    Span4Mux_v I__6576 (
            .O(N__34097),
            .I(N__34082));
    LocalMux I__6575 (
            .O(N__34092),
            .I(N__34082));
    LocalMux I__6574 (
            .O(N__34089),
            .I(N__34082));
    Span4Mux_h I__6573 (
            .O(N__34082),
            .I(N__34079));
    Odrv4 I__6572 (
            .O(N__34079),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__6571 (
            .O(N__34076),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__6570 (
            .O(N__34073),
            .I(N__34070));
    InMux I__6569 (
            .O(N__34070),
            .I(N__34066));
    InMux I__6568 (
            .O(N__34069),
            .I(N__34063));
    LocalMux I__6567 (
            .O(N__34066),
            .I(N__34057));
    LocalMux I__6566 (
            .O(N__34063),
            .I(N__34057));
    InMux I__6565 (
            .O(N__34062),
            .I(N__34054));
    Span4Mux_h I__6564 (
            .O(N__34057),
            .I(N__34051));
    LocalMux I__6563 (
            .O(N__34054),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__6562 (
            .O(N__34051),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__6561 (
            .O(N__34046),
            .I(N__34041));
    InMux I__6560 (
            .O(N__34045),
            .I(N__34038));
    InMux I__6559 (
            .O(N__34044),
            .I(N__34035));
    LocalMux I__6558 (
            .O(N__34041),
            .I(N__34030));
    LocalMux I__6557 (
            .O(N__34038),
            .I(N__34030));
    LocalMux I__6556 (
            .O(N__34035),
            .I(N__34026));
    Span4Mux_v I__6555 (
            .O(N__34030),
            .I(N__34023));
    InMux I__6554 (
            .O(N__34029),
            .I(N__34020));
    Span4Mux_h I__6553 (
            .O(N__34026),
            .I(N__34017));
    Sp12to4 I__6552 (
            .O(N__34023),
            .I(N__34014));
    LocalMux I__6551 (
            .O(N__34020),
            .I(N__34011));
    Odrv4 I__6550 (
            .O(N__34017),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv12 I__6549 (
            .O(N__34014),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv4 I__6548 (
            .O(N__34011),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__6547 (
            .O(N__34004),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__6546 (
            .O(N__34001),
            .I(N__33998));
    InMux I__6545 (
            .O(N__33998),
            .I(N__33994));
    InMux I__6544 (
            .O(N__33997),
            .I(N__33991));
    LocalMux I__6543 (
            .O(N__33994),
            .I(N__33985));
    LocalMux I__6542 (
            .O(N__33991),
            .I(N__33985));
    InMux I__6541 (
            .O(N__33990),
            .I(N__33982));
    Span4Mux_h I__6540 (
            .O(N__33985),
            .I(N__33979));
    LocalMux I__6539 (
            .O(N__33982),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__6538 (
            .O(N__33979),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__6537 (
            .O(N__33974),
            .I(N__33971));
    LocalMux I__6536 (
            .O(N__33971),
            .I(N__33966));
    InMux I__6535 (
            .O(N__33970),
            .I(N__33961));
    InMux I__6534 (
            .O(N__33969),
            .I(N__33961));
    Span4Mux_v I__6533 (
            .O(N__33966),
            .I(N__33955));
    LocalMux I__6532 (
            .O(N__33961),
            .I(N__33955));
    InMux I__6531 (
            .O(N__33960),
            .I(N__33952));
    Span4Mux_h I__6530 (
            .O(N__33955),
            .I(N__33947));
    LocalMux I__6529 (
            .O(N__33952),
            .I(N__33947));
    Sp12to4 I__6528 (
            .O(N__33947),
            .I(N__33944));
    Odrv12 I__6527 (
            .O(N__33944),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__6526 (
            .O(N__33941),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__6525 (
            .O(N__33938),
            .I(N__33935));
    InMux I__6524 (
            .O(N__33935),
            .I(N__33931));
    InMux I__6523 (
            .O(N__33934),
            .I(N__33928));
    LocalMux I__6522 (
            .O(N__33931),
            .I(N__33924));
    LocalMux I__6521 (
            .O(N__33928),
            .I(N__33921));
    InMux I__6520 (
            .O(N__33927),
            .I(N__33918));
    Span4Mux_v I__6519 (
            .O(N__33924),
            .I(N__33915));
    Odrv12 I__6518 (
            .O(N__33921),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__6517 (
            .O(N__33918),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__6516 (
            .O(N__33915),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__6515 (
            .O(N__33908),
            .I(N__33904));
    InMux I__6514 (
            .O(N__33907),
            .I(N__33899));
    LocalMux I__6513 (
            .O(N__33904),
            .I(N__33896));
    InMux I__6512 (
            .O(N__33903),
            .I(N__33891));
    InMux I__6511 (
            .O(N__33902),
            .I(N__33891));
    LocalMux I__6510 (
            .O(N__33899),
            .I(N__33888));
    Span4Mux_v I__6509 (
            .O(N__33896),
            .I(N__33885));
    LocalMux I__6508 (
            .O(N__33891),
            .I(N__33882));
    Span4Mux_h I__6507 (
            .O(N__33888),
            .I(N__33879));
    Sp12to4 I__6506 (
            .O(N__33885),
            .I(N__33874));
    Span12Mux_s9_v I__6505 (
            .O(N__33882),
            .I(N__33874));
    Odrv4 I__6504 (
            .O(N__33879),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv12 I__6503 (
            .O(N__33874),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    CascadeMux I__6502 (
            .O(N__33869),
            .I(N__33866));
    InMux I__6501 (
            .O(N__33866),
            .I(N__33861));
    InMux I__6500 (
            .O(N__33865),
            .I(N__33858));
    InMux I__6499 (
            .O(N__33864),
            .I(N__33855));
    LocalMux I__6498 (
            .O(N__33861),
            .I(N__33852));
    LocalMux I__6497 (
            .O(N__33858),
            .I(N__33849));
    LocalMux I__6496 (
            .O(N__33855),
            .I(N__33844));
    Span4Mux_v I__6495 (
            .O(N__33852),
            .I(N__33844));
    Odrv12 I__6494 (
            .O(N__33849),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__6493 (
            .O(N__33844),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    CascadeMux I__6492 (
            .O(N__33839),
            .I(N__33835));
    InMux I__6491 (
            .O(N__33838),
            .I(N__33831));
    InMux I__6490 (
            .O(N__33835),
            .I(N__33827));
    InMux I__6489 (
            .O(N__33834),
            .I(N__33824));
    LocalMux I__6488 (
            .O(N__33831),
            .I(N__33821));
    InMux I__6487 (
            .O(N__33830),
            .I(N__33818));
    LocalMux I__6486 (
            .O(N__33827),
            .I(N__33815));
    LocalMux I__6485 (
            .O(N__33824),
            .I(N__33808));
    Span4Mux_h I__6484 (
            .O(N__33821),
            .I(N__33808));
    LocalMux I__6483 (
            .O(N__33818),
            .I(N__33808));
    Span4Mux_h I__6482 (
            .O(N__33815),
            .I(N__33805));
    Span4Mux_h I__6481 (
            .O(N__33808),
            .I(N__33802));
    Span4Mux_h I__6480 (
            .O(N__33805),
            .I(N__33799));
    Odrv4 I__6479 (
            .O(N__33802),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv4 I__6478 (
            .O(N__33799),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__6477 (
            .O(N__33794),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__6476 (
            .O(N__33791),
            .I(N__33785));
    InMux I__6475 (
            .O(N__33790),
            .I(N__33785));
    LocalMux I__6474 (
            .O(N__33785),
            .I(N__33781));
    InMux I__6473 (
            .O(N__33784),
            .I(N__33778));
    Span4Mux_h I__6472 (
            .O(N__33781),
            .I(N__33775));
    LocalMux I__6471 (
            .O(N__33778),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__6470 (
            .O(N__33775),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__6469 (
            .O(N__33770),
            .I(N__33765));
    InMux I__6468 (
            .O(N__33769),
            .I(N__33762));
    InMux I__6467 (
            .O(N__33768),
            .I(N__33759));
    LocalMux I__6466 (
            .O(N__33765),
            .I(N__33755));
    LocalMux I__6465 (
            .O(N__33762),
            .I(N__33752));
    LocalMux I__6464 (
            .O(N__33759),
            .I(N__33749));
    InMux I__6463 (
            .O(N__33758),
            .I(N__33746));
    Span4Mux_v I__6462 (
            .O(N__33755),
            .I(N__33743));
    Span4Mux_h I__6461 (
            .O(N__33752),
            .I(N__33740));
    Span4Mux_v I__6460 (
            .O(N__33749),
            .I(N__33737));
    LocalMux I__6459 (
            .O(N__33746),
            .I(N__33734));
    Span4Mux_h I__6458 (
            .O(N__33743),
            .I(N__33729));
    Span4Mux_v I__6457 (
            .O(N__33740),
            .I(N__33729));
    Span4Mux_h I__6456 (
            .O(N__33737),
            .I(N__33724));
    Span4Mux_v I__6455 (
            .O(N__33734),
            .I(N__33724));
    Odrv4 I__6454 (
            .O(N__33729),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__6453 (
            .O(N__33724),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__6452 (
            .O(N__33719),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__6451 (
            .O(N__33716),
            .I(N__33713));
    InMux I__6450 (
            .O(N__33713),
            .I(N__33709));
    InMux I__6449 (
            .O(N__33712),
            .I(N__33706));
    LocalMux I__6448 (
            .O(N__33709),
            .I(N__33700));
    LocalMux I__6447 (
            .O(N__33706),
            .I(N__33700));
    InMux I__6446 (
            .O(N__33705),
            .I(N__33697));
    Span4Mux_h I__6445 (
            .O(N__33700),
            .I(N__33694));
    LocalMux I__6444 (
            .O(N__33697),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__6443 (
            .O(N__33694),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__6442 (
            .O(N__33689),
            .I(N__33684));
    InMux I__6441 (
            .O(N__33688),
            .I(N__33680));
    InMux I__6440 (
            .O(N__33687),
            .I(N__33677));
    LocalMux I__6439 (
            .O(N__33684),
            .I(N__33674));
    InMux I__6438 (
            .O(N__33683),
            .I(N__33671));
    LocalMux I__6437 (
            .O(N__33680),
            .I(N__33666));
    LocalMux I__6436 (
            .O(N__33677),
            .I(N__33666));
    Span4Mux_v I__6435 (
            .O(N__33674),
            .I(N__33663));
    LocalMux I__6434 (
            .O(N__33671),
            .I(N__33660));
    Span4Mux_v I__6433 (
            .O(N__33666),
            .I(N__33657));
    Span4Mux_h I__6432 (
            .O(N__33663),
            .I(N__33652));
    Span4Mux_v I__6431 (
            .O(N__33660),
            .I(N__33652));
    Odrv4 I__6430 (
            .O(N__33657),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__6429 (
            .O(N__33652),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__6428 (
            .O(N__33647),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__6427 (
            .O(N__33644),
            .I(N__33640));
    InMux I__6426 (
            .O(N__33643),
            .I(N__33637));
    InMux I__6425 (
            .O(N__33640),
            .I(N__33634));
    LocalMux I__6424 (
            .O(N__33637),
            .I(N__33628));
    LocalMux I__6423 (
            .O(N__33634),
            .I(N__33628));
    InMux I__6422 (
            .O(N__33633),
            .I(N__33625));
    Span4Mux_h I__6421 (
            .O(N__33628),
            .I(N__33622));
    LocalMux I__6420 (
            .O(N__33625),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv4 I__6419 (
            .O(N__33622),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__6418 (
            .O(N__33617),
            .I(N__33613));
    InMux I__6417 (
            .O(N__33616),
            .I(N__33610));
    LocalMux I__6416 (
            .O(N__33613),
            .I(N__33603));
    LocalMux I__6415 (
            .O(N__33610),
            .I(N__33603));
    InMux I__6414 (
            .O(N__33609),
            .I(N__33600));
    InMux I__6413 (
            .O(N__33608),
            .I(N__33597));
    Span4Mux_v I__6412 (
            .O(N__33603),
            .I(N__33594));
    LocalMux I__6411 (
            .O(N__33600),
            .I(N__33591));
    LocalMux I__6410 (
            .O(N__33597),
            .I(N__33588));
    Span4Mux_h I__6409 (
            .O(N__33594),
            .I(N__33585));
    Span4Mux_v I__6408 (
            .O(N__33591),
            .I(N__33580));
    Span4Mux_v I__6407 (
            .O(N__33588),
            .I(N__33580));
    Odrv4 I__6406 (
            .O(N__33585),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__6405 (
            .O(N__33580),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__6404 (
            .O(N__33575),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__6403 (
            .O(N__33572),
            .I(N__33569));
    InMux I__6402 (
            .O(N__33569),
            .I(N__33565));
    InMux I__6401 (
            .O(N__33568),
            .I(N__33562));
    LocalMux I__6400 (
            .O(N__33565),
            .I(N__33556));
    LocalMux I__6399 (
            .O(N__33562),
            .I(N__33556));
    InMux I__6398 (
            .O(N__33561),
            .I(N__33553));
    Span4Mux_h I__6397 (
            .O(N__33556),
            .I(N__33550));
    LocalMux I__6396 (
            .O(N__33553),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__6395 (
            .O(N__33550),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__6394 (
            .O(N__33545),
            .I(N__33539));
    InMux I__6393 (
            .O(N__33544),
            .I(N__33539));
    LocalMux I__6392 (
            .O(N__33539),
            .I(N__33534));
    InMux I__6391 (
            .O(N__33538),
            .I(N__33531));
    InMux I__6390 (
            .O(N__33537),
            .I(N__33528));
    Span4Mux_h I__6389 (
            .O(N__33534),
            .I(N__33525));
    LocalMux I__6388 (
            .O(N__33531),
            .I(N__33522));
    LocalMux I__6387 (
            .O(N__33528),
            .I(N__33519));
    Span4Mux_h I__6386 (
            .O(N__33525),
            .I(N__33516));
    Span4Mux_h I__6385 (
            .O(N__33522),
            .I(N__33511));
    Span4Mux_h I__6384 (
            .O(N__33519),
            .I(N__33511));
    Odrv4 I__6383 (
            .O(N__33516),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__6382 (
            .O(N__33511),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__6381 (
            .O(N__33506),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__6380 (
            .O(N__33503),
            .I(N__33499));
    CascadeMux I__6379 (
            .O(N__33502),
            .I(N__33496));
    InMux I__6378 (
            .O(N__33499),
            .I(N__33491));
    InMux I__6377 (
            .O(N__33496),
            .I(N__33491));
    LocalMux I__6376 (
            .O(N__33491),
            .I(N__33487));
    InMux I__6375 (
            .O(N__33490),
            .I(N__33484));
    Span4Mux_h I__6374 (
            .O(N__33487),
            .I(N__33481));
    LocalMux I__6373 (
            .O(N__33484),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__6372 (
            .O(N__33481),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__6371 (
            .O(N__33476),
            .I(N__33471));
    InMux I__6370 (
            .O(N__33475),
            .I(N__33466));
    InMux I__6369 (
            .O(N__33474),
            .I(N__33466));
    LocalMux I__6368 (
            .O(N__33471),
            .I(N__33462));
    LocalMux I__6367 (
            .O(N__33466),
            .I(N__33459));
    InMux I__6366 (
            .O(N__33465),
            .I(N__33456));
    Span4Mux_v I__6365 (
            .O(N__33462),
            .I(N__33453));
    Span4Mux_h I__6364 (
            .O(N__33459),
            .I(N__33450));
    LocalMux I__6363 (
            .O(N__33456),
            .I(N__33447));
    Span4Mux_h I__6362 (
            .O(N__33453),
            .I(N__33444));
    Span4Mux_h I__6361 (
            .O(N__33450),
            .I(N__33441));
    Span4Mux_v I__6360 (
            .O(N__33447),
            .I(N__33438));
    Odrv4 I__6359 (
            .O(N__33444),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv4 I__6358 (
            .O(N__33441),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv4 I__6357 (
            .O(N__33438),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__6356 (
            .O(N__33431),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__6355 (
            .O(N__33428),
            .I(N__33425));
    InMux I__6354 (
            .O(N__33425),
            .I(N__33421));
    InMux I__6353 (
            .O(N__33424),
            .I(N__33418));
    LocalMux I__6352 (
            .O(N__33421),
            .I(N__33412));
    LocalMux I__6351 (
            .O(N__33418),
            .I(N__33412));
    InMux I__6350 (
            .O(N__33417),
            .I(N__33409));
    Span4Mux_h I__6349 (
            .O(N__33412),
            .I(N__33406));
    LocalMux I__6348 (
            .O(N__33409),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__6347 (
            .O(N__33406),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    CascadeMux I__6346 (
            .O(N__33401),
            .I(elapsed_time_ns_1_RNIH33T9_0_5_cascade_));
    CascadeMux I__6345 (
            .O(N__33398),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_));
    InMux I__6344 (
            .O(N__33395),
            .I(N__33392));
    LocalMux I__6343 (
            .O(N__33392),
            .I(N__33389));
    Odrv12 I__6342 (
            .O(N__33389),
            .I(\phase_controller_inst1.test_0_sqmuxa ));
    InMux I__6341 (
            .O(N__33386),
            .I(N__33380));
    InMux I__6340 (
            .O(N__33385),
            .I(N__33380));
    LocalMux I__6339 (
            .O(N__33380),
            .I(N__33377));
    Odrv4 I__6338 (
            .O(N__33377),
            .I(\phase_controller_inst1.N_56 ));
    CascadeMux I__6337 (
            .O(N__33374),
            .I(N__33371));
    InMux I__6336 (
            .O(N__33371),
            .I(N__33367));
    InMux I__6335 (
            .O(N__33370),
            .I(N__33364));
    LocalMux I__6334 (
            .O(N__33367),
            .I(N__33360));
    LocalMux I__6333 (
            .O(N__33364),
            .I(N__33357));
    InMux I__6332 (
            .O(N__33363),
            .I(N__33354));
    Span4Mux_h I__6331 (
            .O(N__33360),
            .I(N__33348));
    Span12Mux_h I__6330 (
            .O(N__33357),
            .I(N__33345));
    LocalMux I__6329 (
            .O(N__33354),
            .I(N__33342));
    InMux I__6328 (
            .O(N__33353),
            .I(N__33337));
    InMux I__6327 (
            .O(N__33352),
            .I(N__33337));
    InMux I__6326 (
            .O(N__33351),
            .I(N__33334));
    Span4Mux_v I__6325 (
            .O(N__33348),
            .I(N__33331));
    Span12Mux_v I__6324 (
            .O(N__33345),
            .I(N__33328));
    Span4Mux_h I__6323 (
            .O(N__33342),
            .I(N__33325));
    LocalMux I__6322 (
            .O(N__33337),
            .I(phase_controller_inst1_state_4));
    LocalMux I__6321 (
            .O(N__33334),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__6320 (
            .O(N__33331),
            .I(phase_controller_inst1_state_4));
    Odrv12 I__6319 (
            .O(N__33328),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__6318 (
            .O(N__33325),
            .I(phase_controller_inst1_state_4));
    InMux I__6317 (
            .O(N__33314),
            .I(N__33311));
    LocalMux I__6316 (
            .O(N__33311),
            .I(N__33308));
    Odrv4 I__6315 (
            .O(N__33308),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__6314 (
            .O(N__33305),
            .I(\current_shift_inst.control_input_cry_24 ));
    CascadeMux I__6313 (
            .O(N__33302),
            .I(N__33299));
    InMux I__6312 (
            .O(N__33299),
            .I(N__33296));
    LocalMux I__6311 (
            .O(N__33296),
            .I(N__33293));
    Odrv4 I__6310 (
            .O(N__33293),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ));
    InMux I__6309 (
            .O(N__33290),
            .I(\current_shift_inst.control_input_cry_25 ));
    InMux I__6308 (
            .O(N__33287),
            .I(N__33284));
    LocalMux I__6307 (
            .O(N__33284),
            .I(N__33281));
    Odrv4 I__6306 (
            .O(N__33281),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ));
    InMux I__6305 (
            .O(N__33278),
            .I(\current_shift_inst.control_input_cry_26 ));
    InMux I__6304 (
            .O(N__33275),
            .I(N__33272));
    LocalMux I__6303 (
            .O(N__33272),
            .I(N__33269));
    Odrv4 I__6302 (
            .O(N__33269),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ));
    InMux I__6301 (
            .O(N__33266),
            .I(\current_shift_inst.control_input_cry_27 ));
    CascadeMux I__6300 (
            .O(N__33263),
            .I(N__33260));
    InMux I__6299 (
            .O(N__33260),
            .I(N__33257));
    LocalMux I__6298 (
            .O(N__33257),
            .I(N__33254));
    Odrv4 I__6297 (
            .O(N__33254),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ));
    InMux I__6296 (
            .O(N__33251),
            .I(\current_shift_inst.control_input_cry_28 ));
    InMux I__6295 (
            .O(N__33248),
            .I(\current_shift_inst.control_input_cry_29 ));
    InMux I__6294 (
            .O(N__33245),
            .I(N__33242));
    LocalMux I__6293 (
            .O(N__33242),
            .I(N__33238));
    InMux I__6292 (
            .O(N__33241),
            .I(N__33235));
    Odrv4 I__6291 (
            .O(N__33238),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__6290 (
            .O(N__33235),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__6289 (
            .O(N__33230),
            .I(N__33227));
    LocalMux I__6288 (
            .O(N__33227),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ));
    IoInMux I__6287 (
            .O(N__33224),
            .I(N__33221));
    LocalMux I__6286 (
            .O(N__33221),
            .I(N__33218));
    Span4Mux_s0_v I__6285 (
            .O(N__33218),
            .I(N__33215));
    Odrv4 I__6284 (
            .O(N__33215),
            .I(\pll_inst.red_c_i ));
    InMux I__6283 (
            .O(N__33212),
            .I(N__33208));
    InMux I__6282 (
            .O(N__33211),
            .I(N__33204));
    LocalMux I__6281 (
            .O(N__33208),
            .I(N__33201));
    InMux I__6280 (
            .O(N__33207),
            .I(N__33198));
    LocalMux I__6279 (
            .O(N__33204),
            .I(N__33195));
    Span4Mux_v I__6278 (
            .O(N__33201),
            .I(N__33190));
    LocalMux I__6277 (
            .O(N__33198),
            .I(N__33190));
    Span12Mux_h I__6276 (
            .O(N__33195),
            .I(N__33187));
    Span4Mux_h I__6275 (
            .O(N__33190),
            .I(N__33184));
    Span12Mux_v I__6274 (
            .O(N__33187),
            .I(N__33181));
    Span4Mux_v I__6273 (
            .O(N__33184),
            .I(N__33178));
    Odrv12 I__6272 (
            .O(N__33181),
            .I(il_min_comp1_c));
    Odrv4 I__6271 (
            .O(N__33178),
            .I(il_min_comp1_c));
    InMux I__6270 (
            .O(N__33173),
            .I(N__33170));
    LocalMux I__6269 (
            .O(N__33170),
            .I(N__33167));
    Odrv4 I__6268 (
            .O(N__33167),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__6267 (
            .O(N__33164),
            .I(\current_shift_inst.control_input_cry_16 ));
    CascadeMux I__6266 (
            .O(N__33161),
            .I(N__33158));
    InMux I__6265 (
            .O(N__33158),
            .I(N__33155));
    LocalMux I__6264 (
            .O(N__33155),
            .I(N__33152));
    Odrv4 I__6263 (
            .O(N__33152),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    InMux I__6262 (
            .O(N__33149),
            .I(\current_shift_inst.control_input_cry_17 ));
    InMux I__6261 (
            .O(N__33146),
            .I(N__33143));
    LocalMux I__6260 (
            .O(N__33143),
            .I(N__33140));
    Odrv4 I__6259 (
            .O(N__33140),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__6258 (
            .O(N__33137),
            .I(\current_shift_inst.control_input_cry_18 ));
    InMux I__6257 (
            .O(N__33134),
            .I(N__33131));
    LocalMux I__6256 (
            .O(N__33131),
            .I(N__33128));
    Odrv4 I__6255 (
            .O(N__33128),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__6254 (
            .O(N__33125),
            .I(\current_shift_inst.control_input_cry_19 ));
    CascadeMux I__6253 (
            .O(N__33122),
            .I(N__33119));
    InMux I__6252 (
            .O(N__33119),
            .I(N__33116));
    LocalMux I__6251 (
            .O(N__33116),
            .I(N__33113));
    Odrv4 I__6250 (
            .O(N__33113),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__6249 (
            .O(N__33110),
            .I(\current_shift_inst.control_input_cry_20 ));
    InMux I__6248 (
            .O(N__33107),
            .I(N__33104));
    LocalMux I__6247 (
            .O(N__33104),
            .I(N__33101));
    Odrv4 I__6246 (
            .O(N__33101),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__6245 (
            .O(N__33098),
            .I(\current_shift_inst.control_input_cry_21 ));
    CascadeMux I__6244 (
            .O(N__33095),
            .I(N__33092));
    InMux I__6243 (
            .O(N__33092),
            .I(N__33089));
    LocalMux I__6242 (
            .O(N__33089),
            .I(N__33086));
    Odrv4 I__6241 (
            .O(N__33086),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__6240 (
            .O(N__33083),
            .I(\current_shift_inst.control_input_cry_22 ));
    CascadeMux I__6239 (
            .O(N__33080),
            .I(N__33077));
    InMux I__6238 (
            .O(N__33077),
            .I(N__33074));
    LocalMux I__6237 (
            .O(N__33074),
            .I(N__33071));
    Odrv4 I__6236 (
            .O(N__33071),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__6235 (
            .O(N__33068),
            .I(bfn_12_20_0_));
    CascadeMux I__6234 (
            .O(N__33065),
            .I(N__33062));
    InMux I__6233 (
            .O(N__33062),
            .I(N__33059));
    LocalMux I__6232 (
            .O(N__33059),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__6231 (
            .O(N__33056),
            .I(N__33053));
    LocalMux I__6230 (
            .O(N__33053),
            .I(N__33050));
    Odrv4 I__6229 (
            .O(N__33050),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__6228 (
            .O(N__33047),
            .I(\current_shift_inst.control_input_cry_8 ));
    CascadeMux I__6227 (
            .O(N__33044),
            .I(N__33041));
    InMux I__6226 (
            .O(N__33041),
            .I(N__33038));
    LocalMux I__6225 (
            .O(N__33038),
            .I(N__33035));
    Odrv4 I__6224 (
            .O(N__33035),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__6223 (
            .O(N__33032),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__6222 (
            .O(N__33029),
            .I(N__33026));
    LocalMux I__6221 (
            .O(N__33026),
            .I(N__33023));
    Odrv4 I__6220 (
            .O(N__33023),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__6219 (
            .O(N__33020),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__6218 (
            .O(N__33017),
            .I(N__33014));
    LocalMux I__6217 (
            .O(N__33014),
            .I(N__33011));
    Odrv4 I__6216 (
            .O(N__33011),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__6215 (
            .O(N__33008),
            .I(\current_shift_inst.control_input_cry_11 ));
    CascadeMux I__6214 (
            .O(N__33005),
            .I(N__33002));
    InMux I__6213 (
            .O(N__33002),
            .I(N__32999));
    LocalMux I__6212 (
            .O(N__32999),
            .I(N__32996));
    Odrv4 I__6211 (
            .O(N__32996),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__6210 (
            .O(N__32993),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__6209 (
            .O(N__32990),
            .I(N__32987));
    LocalMux I__6208 (
            .O(N__32987),
            .I(N__32984));
    Odrv4 I__6207 (
            .O(N__32984),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__6206 (
            .O(N__32981),
            .I(\current_shift_inst.control_input_cry_13 ));
    CascadeMux I__6205 (
            .O(N__32978),
            .I(N__32975));
    InMux I__6204 (
            .O(N__32975),
            .I(N__32972));
    LocalMux I__6203 (
            .O(N__32972),
            .I(N__32969));
    Odrv4 I__6202 (
            .O(N__32969),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__6201 (
            .O(N__32966),
            .I(\current_shift_inst.control_input_cry_14 ));
    CascadeMux I__6200 (
            .O(N__32963),
            .I(N__32960));
    InMux I__6199 (
            .O(N__32960),
            .I(N__32957));
    LocalMux I__6198 (
            .O(N__32957),
            .I(N__32954));
    Odrv4 I__6197 (
            .O(N__32954),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__6196 (
            .O(N__32951),
            .I(bfn_12_19_0_));
    InMux I__6195 (
            .O(N__32948),
            .I(N__32945));
    LocalMux I__6194 (
            .O(N__32945),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__6193 (
            .O(N__32942),
            .I(N__32939));
    InMux I__6192 (
            .O(N__32939),
            .I(N__32936));
    LocalMux I__6191 (
            .O(N__32936),
            .I(N__32931));
    InMux I__6190 (
            .O(N__32935),
            .I(N__32928));
    InMux I__6189 (
            .O(N__32934),
            .I(N__32925));
    Span4Mux_h I__6188 (
            .O(N__32931),
            .I(N__32922));
    LocalMux I__6187 (
            .O(N__32928),
            .I(\current_shift_inst.N_1271_i ));
    LocalMux I__6186 (
            .O(N__32925),
            .I(\current_shift_inst.N_1271_i ));
    Odrv4 I__6185 (
            .O(N__32922),
            .I(\current_shift_inst.N_1271_i ));
    InMux I__6184 (
            .O(N__32915),
            .I(N__32912));
    LocalMux I__6183 (
            .O(N__32912),
            .I(N__32909));
    Odrv4 I__6182 (
            .O(N__32909),
            .I(\current_shift_inst.control_input_1 ));
    InMux I__6181 (
            .O(N__32906),
            .I(N__32903));
    LocalMux I__6180 (
            .O(N__32903),
            .I(N__32900));
    Odrv4 I__6179 (
            .O(N__32900),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__6178 (
            .O(N__32897),
            .I(\current_shift_inst.control_input_cry_0 ));
    CascadeMux I__6177 (
            .O(N__32894),
            .I(N__32891));
    InMux I__6176 (
            .O(N__32891),
            .I(N__32888));
    LocalMux I__6175 (
            .O(N__32888),
            .I(N__32885));
    Odrv4 I__6174 (
            .O(N__32885),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__6173 (
            .O(N__32882),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__6172 (
            .O(N__32879),
            .I(N__32876));
    LocalMux I__6171 (
            .O(N__32876),
            .I(N__32873));
    Odrv4 I__6170 (
            .O(N__32873),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__6169 (
            .O(N__32870),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__6168 (
            .O(N__32867),
            .I(N__32864));
    LocalMux I__6167 (
            .O(N__32864),
            .I(N__32861));
    Odrv4 I__6166 (
            .O(N__32861),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__6165 (
            .O(N__32858),
            .I(\current_shift_inst.control_input_cry_3 ));
    CascadeMux I__6164 (
            .O(N__32855),
            .I(N__32852));
    InMux I__6163 (
            .O(N__32852),
            .I(N__32849));
    LocalMux I__6162 (
            .O(N__32849),
            .I(N__32846));
    Odrv4 I__6161 (
            .O(N__32846),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__6160 (
            .O(N__32843),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__6159 (
            .O(N__32840),
            .I(N__32837));
    LocalMux I__6158 (
            .O(N__32837),
            .I(N__32834));
    Odrv4 I__6157 (
            .O(N__32834),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__6156 (
            .O(N__32831),
            .I(\current_shift_inst.control_input_cry_5 ));
    CascadeMux I__6155 (
            .O(N__32828),
            .I(N__32825));
    InMux I__6154 (
            .O(N__32825),
            .I(N__32822));
    LocalMux I__6153 (
            .O(N__32822),
            .I(N__32819));
    Odrv4 I__6152 (
            .O(N__32819),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__6151 (
            .O(N__32816),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__6150 (
            .O(N__32813),
            .I(N__32810));
    LocalMux I__6149 (
            .O(N__32810),
            .I(\current_shift_inst.control_input_axb_8 ));
    CascadeMux I__6148 (
            .O(N__32807),
            .I(N__32804));
    InMux I__6147 (
            .O(N__32804),
            .I(N__32801));
    LocalMux I__6146 (
            .O(N__32801),
            .I(N__32798));
    Odrv4 I__6145 (
            .O(N__32798),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__6144 (
            .O(N__32795),
            .I(bfn_12_18_0_));
    InMux I__6143 (
            .O(N__32792),
            .I(N__32785));
    InMux I__6142 (
            .O(N__32791),
            .I(N__32785));
    InMux I__6141 (
            .O(N__32790),
            .I(N__32782));
    LocalMux I__6140 (
            .O(N__32785),
            .I(N__32779));
    LocalMux I__6139 (
            .O(N__32782),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__6138 (
            .O(N__32779),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__6137 (
            .O(N__32774),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    CascadeMux I__6136 (
            .O(N__32771),
            .I(N__32767));
    CascadeMux I__6135 (
            .O(N__32770),
            .I(N__32764));
    InMux I__6134 (
            .O(N__32767),
            .I(N__32761));
    InMux I__6133 (
            .O(N__32764),
            .I(N__32757));
    LocalMux I__6132 (
            .O(N__32761),
            .I(N__32754));
    InMux I__6131 (
            .O(N__32760),
            .I(N__32751));
    LocalMux I__6130 (
            .O(N__32757),
            .I(N__32746));
    Span4Mux_h I__6129 (
            .O(N__32754),
            .I(N__32746));
    LocalMux I__6128 (
            .O(N__32751),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__6127 (
            .O(N__32746),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__6126 (
            .O(N__32741),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    CEMux I__6125 (
            .O(N__32738),
            .I(N__32733));
    CEMux I__6124 (
            .O(N__32737),
            .I(N__32730));
    CEMux I__6123 (
            .O(N__32736),
            .I(N__32727));
    LocalMux I__6122 (
            .O(N__32733),
            .I(N__32716));
    LocalMux I__6121 (
            .O(N__32730),
            .I(N__32716));
    LocalMux I__6120 (
            .O(N__32727),
            .I(N__32699));
    CEMux I__6119 (
            .O(N__32726),
            .I(N__32696));
    CEMux I__6118 (
            .O(N__32725),
            .I(N__32693));
    InMux I__6117 (
            .O(N__32724),
            .I(N__32680));
    InMux I__6116 (
            .O(N__32723),
            .I(N__32680));
    InMux I__6115 (
            .O(N__32722),
            .I(N__32680));
    CEMux I__6114 (
            .O(N__32721),
            .I(N__32676));
    Span4Mux_v I__6113 (
            .O(N__32716),
            .I(N__32662));
    InMux I__6112 (
            .O(N__32715),
            .I(N__32653));
    InMux I__6111 (
            .O(N__32714),
            .I(N__32653));
    InMux I__6110 (
            .O(N__32713),
            .I(N__32653));
    InMux I__6109 (
            .O(N__32712),
            .I(N__32653));
    InMux I__6108 (
            .O(N__32711),
            .I(N__32644));
    InMux I__6107 (
            .O(N__32710),
            .I(N__32644));
    InMux I__6106 (
            .O(N__32709),
            .I(N__32644));
    InMux I__6105 (
            .O(N__32708),
            .I(N__32644));
    InMux I__6104 (
            .O(N__32707),
            .I(N__32635));
    InMux I__6103 (
            .O(N__32706),
            .I(N__32635));
    InMux I__6102 (
            .O(N__32705),
            .I(N__32635));
    InMux I__6101 (
            .O(N__32704),
            .I(N__32635));
    CEMux I__6100 (
            .O(N__32703),
            .I(N__32632));
    CEMux I__6099 (
            .O(N__32702),
            .I(N__32628));
    Span4Mux_v I__6098 (
            .O(N__32699),
            .I(N__32620));
    LocalMux I__6097 (
            .O(N__32696),
            .I(N__32620));
    LocalMux I__6096 (
            .O(N__32693),
            .I(N__32620));
    InMux I__6095 (
            .O(N__32692),
            .I(N__32611));
    InMux I__6094 (
            .O(N__32691),
            .I(N__32611));
    InMux I__6093 (
            .O(N__32690),
            .I(N__32611));
    InMux I__6092 (
            .O(N__32689),
            .I(N__32611));
    InMux I__6091 (
            .O(N__32688),
            .I(N__32608));
    CEMux I__6090 (
            .O(N__32687),
            .I(N__32605));
    LocalMux I__6089 (
            .O(N__32680),
            .I(N__32602));
    CEMux I__6088 (
            .O(N__32679),
            .I(N__32599));
    LocalMux I__6087 (
            .O(N__32676),
            .I(N__32596));
    InMux I__6086 (
            .O(N__32675),
            .I(N__32587));
    InMux I__6085 (
            .O(N__32674),
            .I(N__32587));
    InMux I__6084 (
            .O(N__32673),
            .I(N__32587));
    InMux I__6083 (
            .O(N__32672),
            .I(N__32587));
    InMux I__6082 (
            .O(N__32671),
            .I(N__32580));
    InMux I__6081 (
            .O(N__32670),
            .I(N__32580));
    InMux I__6080 (
            .O(N__32669),
            .I(N__32580));
    InMux I__6079 (
            .O(N__32668),
            .I(N__32571));
    InMux I__6078 (
            .O(N__32667),
            .I(N__32571));
    InMux I__6077 (
            .O(N__32666),
            .I(N__32571));
    InMux I__6076 (
            .O(N__32665),
            .I(N__32571));
    Span4Mux_v I__6075 (
            .O(N__32662),
            .I(N__32564));
    LocalMux I__6074 (
            .O(N__32653),
            .I(N__32564));
    LocalMux I__6073 (
            .O(N__32644),
            .I(N__32564));
    LocalMux I__6072 (
            .O(N__32635),
            .I(N__32561));
    LocalMux I__6071 (
            .O(N__32632),
            .I(N__32557));
    CEMux I__6070 (
            .O(N__32631),
            .I(N__32554));
    LocalMux I__6069 (
            .O(N__32628),
            .I(N__32551));
    CEMux I__6068 (
            .O(N__32627),
            .I(N__32548));
    Span4Mux_h I__6067 (
            .O(N__32620),
            .I(N__32545));
    LocalMux I__6066 (
            .O(N__32611),
            .I(N__32542));
    LocalMux I__6065 (
            .O(N__32608),
            .I(N__32539));
    LocalMux I__6064 (
            .O(N__32605),
            .I(N__32534));
    Span4Mux_h I__6063 (
            .O(N__32602),
            .I(N__32534));
    LocalMux I__6062 (
            .O(N__32599),
            .I(N__32529));
    Span4Mux_v I__6061 (
            .O(N__32596),
            .I(N__32529));
    LocalMux I__6060 (
            .O(N__32587),
            .I(N__32518));
    LocalMux I__6059 (
            .O(N__32580),
            .I(N__32518));
    LocalMux I__6058 (
            .O(N__32571),
            .I(N__32518));
    Span4Mux_h I__6057 (
            .O(N__32564),
            .I(N__32518));
    Span4Mux_v I__6056 (
            .O(N__32561),
            .I(N__32518));
    CEMux I__6055 (
            .O(N__32560),
            .I(N__32515));
    Span4Mux_v I__6054 (
            .O(N__32557),
            .I(N__32512));
    LocalMux I__6053 (
            .O(N__32554),
            .I(N__32507));
    Sp12to4 I__6052 (
            .O(N__32551),
            .I(N__32507));
    LocalMux I__6051 (
            .O(N__32548),
            .I(N__32500));
    Span4Mux_v I__6050 (
            .O(N__32545),
            .I(N__32500));
    Span4Mux_h I__6049 (
            .O(N__32542),
            .I(N__32500));
    Span4Mux_h I__6048 (
            .O(N__32539),
            .I(N__32495));
    Span4Mux_v I__6047 (
            .O(N__32534),
            .I(N__32495));
    Span4Mux_v I__6046 (
            .O(N__32529),
            .I(N__32490));
    Span4Mux_v I__6045 (
            .O(N__32518),
            .I(N__32490));
    LocalMux I__6044 (
            .O(N__32515),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6043 (
            .O(N__32512),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv12 I__6042 (
            .O(N__32507),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6041 (
            .O(N__32500),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6040 (
            .O(N__32495),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__6039 (
            .O(N__32490),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__6038 (
            .O(N__32477),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__6037 (
            .O(N__32474),
            .I(N__32469));
    InMux I__6036 (
            .O(N__32473),
            .I(N__32466));
    InMux I__6035 (
            .O(N__32472),
            .I(N__32463));
    LocalMux I__6034 (
            .O(N__32469),
            .I(N__32458));
    LocalMux I__6033 (
            .O(N__32466),
            .I(N__32458));
    LocalMux I__6032 (
            .O(N__32463),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv12 I__6031 (
            .O(N__32458),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__6030 (
            .O(N__32453),
            .I(N__32450));
    LocalMux I__6029 (
            .O(N__32450),
            .I(N__32445));
    InMux I__6028 (
            .O(N__32449),
            .I(N__32442));
    InMux I__6027 (
            .O(N__32448),
            .I(N__32439));
    Span4Mux_h I__6026 (
            .O(N__32445),
            .I(N__32436));
    LocalMux I__6025 (
            .O(N__32442),
            .I(N__32433));
    LocalMux I__6024 (
            .O(N__32439),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    Odrv4 I__6023 (
            .O(N__32436),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    Odrv12 I__6022 (
            .O(N__32433),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__6021 (
            .O(N__32426),
            .I(N__32387));
    InMux I__6020 (
            .O(N__32425),
            .I(N__32387));
    InMux I__6019 (
            .O(N__32424),
            .I(N__32380));
    InMux I__6018 (
            .O(N__32423),
            .I(N__32380));
    InMux I__6017 (
            .O(N__32422),
            .I(N__32380));
    InMux I__6016 (
            .O(N__32421),
            .I(N__32373));
    InMux I__6015 (
            .O(N__32420),
            .I(N__32373));
    InMux I__6014 (
            .O(N__32419),
            .I(N__32373));
    InMux I__6013 (
            .O(N__32418),
            .I(N__32368));
    InMux I__6012 (
            .O(N__32417),
            .I(N__32368));
    InMux I__6011 (
            .O(N__32416),
            .I(N__32363));
    InMux I__6010 (
            .O(N__32415),
            .I(N__32363));
    InMux I__6009 (
            .O(N__32414),
            .I(N__32341));
    InMux I__6008 (
            .O(N__32413),
            .I(N__32319));
    InMux I__6007 (
            .O(N__32412),
            .I(N__32319));
    InMux I__6006 (
            .O(N__32411),
            .I(N__32316));
    InMux I__6005 (
            .O(N__32410),
            .I(N__32313));
    InMux I__6004 (
            .O(N__32409),
            .I(N__32310));
    InMux I__6003 (
            .O(N__32408),
            .I(N__32300));
    InMux I__6002 (
            .O(N__32407),
            .I(N__32291));
    InMux I__6001 (
            .O(N__32406),
            .I(N__32291));
    InMux I__6000 (
            .O(N__32405),
            .I(N__32291));
    InMux I__5999 (
            .O(N__32404),
            .I(N__32291));
    InMux I__5998 (
            .O(N__32403),
            .I(N__32278));
    InMux I__5997 (
            .O(N__32402),
            .I(N__32278));
    InMux I__5996 (
            .O(N__32401),
            .I(N__32278));
    InMux I__5995 (
            .O(N__32400),
            .I(N__32278));
    InMux I__5994 (
            .O(N__32399),
            .I(N__32278));
    InMux I__5993 (
            .O(N__32398),
            .I(N__32278));
    InMux I__5992 (
            .O(N__32397),
            .I(N__32269));
    InMux I__5991 (
            .O(N__32396),
            .I(N__32269));
    InMux I__5990 (
            .O(N__32395),
            .I(N__32269));
    InMux I__5989 (
            .O(N__32394),
            .I(N__32269));
    InMux I__5988 (
            .O(N__32393),
            .I(N__32264));
    InMux I__5987 (
            .O(N__32392),
            .I(N__32264));
    LocalMux I__5986 (
            .O(N__32387),
            .I(N__32253));
    LocalMux I__5985 (
            .O(N__32380),
            .I(N__32253));
    LocalMux I__5984 (
            .O(N__32373),
            .I(N__32253));
    LocalMux I__5983 (
            .O(N__32368),
            .I(N__32253));
    LocalMux I__5982 (
            .O(N__32363),
            .I(N__32253));
    InMux I__5981 (
            .O(N__32362),
            .I(N__32242));
    InMux I__5980 (
            .O(N__32361),
            .I(N__32242));
    InMux I__5979 (
            .O(N__32360),
            .I(N__32242));
    InMux I__5978 (
            .O(N__32359),
            .I(N__32242));
    InMux I__5977 (
            .O(N__32358),
            .I(N__32242));
    InMux I__5976 (
            .O(N__32357),
            .I(N__32239));
    InMux I__5975 (
            .O(N__32356),
            .I(N__32228));
    InMux I__5974 (
            .O(N__32355),
            .I(N__32228));
    InMux I__5973 (
            .O(N__32354),
            .I(N__32228));
    InMux I__5972 (
            .O(N__32353),
            .I(N__32228));
    InMux I__5971 (
            .O(N__32352),
            .I(N__32228));
    InMux I__5970 (
            .O(N__32351),
            .I(N__32217));
    InMux I__5969 (
            .O(N__32350),
            .I(N__32217));
    InMux I__5968 (
            .O(N__32349),
            .I(N__32217));
    InMux I__5967 (
            .O(N__32348),
            .I(N__32217));
    InMux I__5966 (
            .O(N__32347),
            .I(N__32217));
    InMux I__5965 (
            .O(N__32346),
            .I(N__32210));
    InMux I__5964 (
            .O(N__32345),
            .I(N__32210));
    InMux I__5963 (
            .O(N__32344),
            .I(N__32210));
    LocalMux I__5962 (
            .O(N__32341),
            .I(N__32207));
    InMux I__5961 (
            .O(N__32340),
            .I(N__32200));
    InMux I__5960 (
            .O(N__32339),
            .I(N__32200));
    InMux I__5959 (
            .O(N__32338),
            .I(N__32200));
    InMux I__5958 (
            .O(N__32337),
            .I(N__32191));
    InMux I__5957 (
            .O(N__32336),
            .I(N__32191));
    InMux I__5956 (
            .O(N__32335),
            .I(N__32191));
    InMux I__5955 (
            .O(N__32334),
            .I(N__32191));
    InMux I__5954 (
            .O(N__32333),
            .I(N__32171));
    InMux I__5953 (
            .O(N__32332),
            .I(N__32171));
    InMux I__5952 (
            .O(N__32331),
            .I(N__32171));
    InMux I__5951 (
            .O(N__32330),
            .I(N__32171));
    InMux I__5950 (
            .O(N__32329),
            .I(N__32171));
    InMux I__5949 (
            .O(N__32328),
            .I(N__32171));
    InMux I__5948 (
            .O(N__32327),
            .I(N__32161));
    InMux I__5947 (
            .O(N__32326),
            .I(N__32156));
    InMux I__5946 (
            .O(N__32325),
            .I(N__32156));
    InMux I__5945 (
            .O(N__32324),
            .I(N__32153));
    LocalMux I__5944 (
            .O(N__32319),
            .I(N__32150));
    LocalMux I__5943 (
            .O(N__32316),
            .I(N__32143));
    LocalMux I__5942 (
            .O(N__32313),
            .I(N__32143));
    LocalMux I__5941 (
            .O(N__32310),
            .I(N__32143));
    InMux I__5940 (
            .O(N__32309),
            .I(N__32128));
    InMux I__5939 (
            .O(N__32308),
            .I(N__32128));
    InMux I__5938 (
            .O(N__32307),
            .I(N__32128));
    InMux I__5937 (
            .O(N__32306),
            .I(N__32128));
    InMux I__5936 (
            .O(N__32305),
            .I(N__32128));
    InMux I__5935 (
            .O(N__32304),
            .I(N__32128));
    InMux I__5934 (
            .O(N__32303),
            .I(N__32128));
    LocalMux I__5933 (
            .O(N__32300),
            .I(N__32115));
    LocalMux I__5932 (
            .O(N__32291),
            .I(N__32115));
    LocalMux I__5931 (
            .O(N__32278),
            .I(N__32115));
    LocalMux I__5930 (
            .O(N__32269),
            .I(N__32115));
    LocalMux I__5929 (
            .O(N__32264),
            .I(N__32115));
    Span4Mux_v I__5928 (
            .O(N__32253),
            .I(N__32115));
    LocalMux I__5927 (
            .O(N__32242),
            .I(N__32112));
    LocalMux I__5926 (
            .O(N__32239),
            .I(N__32107));
    LocalMux I__5925 (
            .O(N__32228),
            .I(N__32107));
    LocalMux I__5924 (
            .O(N__32217),
            .I(N__32096));
    LocalMux I__5923 (
            .O(N__32210),
            .I(N__32096));
    Span4Mux_v I__5922 (
            .O(N__32207),
            .I(N__32096));
    LocalMux I__5921 (
            .O(N__32200),
            .I(N__32096));
    LocalMux I__5920 (
            .O(N__32191),
            .I(N__32096));
    InMux I__5919 (
            .O(N__32190),
            .I(N__32093));
    InMux I__5918 (
            .O(N__32189),
            .I(N__32090));
    InMux I__5917 (
            .O(N__32188),
            .I(N__32079));
    InMux I__5916 (
            .O(N__32187),
            .I(N__32079));
    InMux I__5915 (
            .O(N__32186),
            .I(N__32079));
    InMux I__5914 (
            .O(N__32185),
            .I(N__32079));
    InMux I__5913 (
            .O(N__32184),
            .I(N__32079));
    LocalMux I__5912 (
            .O(N__32171),
            .I(N__32076));
    InMux I__5911 (
            .O(N__32170),
            .I(N__32067));
    InMux I__5910 (
            .O(N__32169),
            .I(N__32067));
    InMux I__5909 (
            .O(N__32168),
            .I(N__32067));
    InMux I__5908 (
            .O(N__32167),
            .I(N__32067));
    InMux I__5907 (
            .O(N__32166),
            .I(N__32062));
    InMux I__5906 (
            .O(N__32165),
            .I(N__32062));
    InMux I__5905 (
            .O(N__32164),
            .I(N__32059));
    LocalMux I__5904 (
            .O(N__32161),
            .I(N__32054));
    LocalMux I__5903 (
            .O(N__32156),
            .I(N__32054));
    LocalMux I__5902 (
            .O(N__32153),
            .I(N__32051));
    Span4Mux_v I__5901 (
            .O(N__32150),
            .I(N__32048));
    Span4Mux_v I__5900 (
            .O(N__32143),
            .I(N__32041));
    LocalMux I__5899 (
            .O(N__32128),
            .I(N__32041));
    Span4Mux_v I__5898 (
            .O(N__32115),
            .I(N__32041));
    Span12Mux_s11_h I__5897 (
            .O(N__32112),
            .I(N__32038));
    Span4Mux_h I__5896 (
            .O(N__32107),
            .I(N__32033));
    Span4Mux_v I__5895 (
            .O(N__32096),
            .I(N__32033));
    LocalMux I__5894 (
            .O(N__32093),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5893 (
            .O(N__32090),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5892 (
            .O(N__32079),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5891 (
            .O(N__32076),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5890 (
            .O(N__32067),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5889 (
            .O(N__32062),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5888 (
            .O(N__32059),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5887 (
            .O(N__32054),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5886 (
            .O(N__32051),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5885 (
            .O(N__32048),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5884 (
            .O(N__32041),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__5883 (
            .O(N__32038),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5882 (
            .O(N__32033),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__5881 (
            .O(N__32006),
            .I(N__32003));
    LocalMux I__5880 (
            .O(N__32003),
            .I(N__31998));
    InMux I__5879 (
            .O(N__32002),
            .I(N__31995));
    InMux I__5878 (
            .O(N__32001),
            .I(N__31992));
    Span4Mux_h I__5877 (
            .O(N__31998),
            .I(N__31989));
    LocalMux I__5876 (
            .O(N__31995),
            .I(N__31986));
    LocalMux I__5875 (
            .O(N__31992),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    Odrv4 I__5874 (
            .O(N__31989),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    Odrv4 I__5873 (
            .O(N__31986),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    InMux I__5872 (
            .O(N__31979),
            .I(N__31976));
    LocalMux I__5871 (
            .O(N__31976),
            .I(N__31972));
    InMux I__5870 (
            .O(N__31975),
            .I(N__31969));
    Odrv12 I__5869 (
            .O(N__31972),
            .I(\phase_controller_inst1.N_52 ));
    LocalMux I__5868 (
            .O(N__31969),
            .I(\phase_controller_inst1.N_52 ));
    InMux I__5867 (
            .O(N__31964),
            .I(N__31961));
    LocalMux I__5866 (
            .O(N__31961),
            .I(phase_controller_inst1_N_54));
    CascadeMux I__5865 (
            .O(N__31958),
            .I(N__31955));
    InMux I__5864 (
            .O(N__31955),
            .I(N__31951));
    InMux I__5863 (
            .O(N__31954),
            .I(N__31947));
    LocalMux I__5862 (
            .O(N__31951),
            .I(N__31942));
    InMux I__5861 (
            .O(N__31950),
            .I(N__31939));
    LocalMux I__5860 (
            .O(N__31947),
            .I(N__31936));
    InMux I__5859 (
            .O(N__31946),
            .I(N__31933));
    InMux I__5858 (
            .O(N__31945),
            .I(N__31930));
    Span4Mux_v I__5857 (
            .O(N__31942),
            .I(N__31925));
    LocalMux I__5856 (
            .O(N__31939),
            .I(N__31925));
    Span4Mux_v I__5855 (
            .O(N__31936),
            .I(N__31922));
    LocalMux I__5854 (
            .O(N__31933),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__5853 (
            .O(N__31930),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__5852 (
            .O(N__31925),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__5851 (
            .O(N__31922),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    InMux I__5850 (
            .O(N__31913),
            .I(N__31909));
    InMux I__5849 (
            .O(N__31912),
            .I(N__31906));
    LocalMux I__5848 (
            .O(N__31909),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    LocalMux I__5847 (
            .O(N__31906),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__5846 (
            .O(N__31901),
            .I(N__31897));
    InMux I__5845 (
            .O(N__31900),
            .I(N__31893));
    LocalMux I__5844 (
            .O(N__31897),
            .I(N__31890));
    InMux I__5843 (
            .O(N__31896),
            .I(N__31887));
    LocalMux I__5842 (
            .O(N__31893),
            .I(N__31884));
    Span4Mux_h I__5841 (
            .O(N__31890),
            .I(N__31881));
    LocalMux I__5840 (
            .O(N__31887),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__5839 (
            .O(N__31884),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__5838 (
            .O(N__31881),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__5837 (
            .O(N__31874),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__5836 (
            .O(N__31871),
            .I(N__31867));
    InMux I__5835 (
            .O(N__31870),
            .I(N__31863));
    LocalMux I__5834 (
            .O(N__31867),
            .I(N__31860));
    InMux I__5833 (
            .O(N__31866),
            .I(N__31857));
    LocalMux I__5832 (
            .O(N__31863),
            .I(N__31852));
    Span4Mux_v I__5831 (
            .O(N__31860),
            .I(N__31852));
    LocalMux I__5830 (
            .O(N__31857),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__5829 (
            .O(N__31852),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__5828 (
            .O(N__31847),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__5827 (
            .O(N__31844),
            .I(N__31838));
    InMux I__5826 (
            .O(N__31843),
            .I(N__31838));
    LocalMux I__5825 (
            .O(N__31838),
            .I(N__31834));
    InMux I__5824 (
            .O(N__31837),
            .I(N__31831));
    Span4Mux_h I__5823 (
            .O(N__31834),
            .I(N__31828));
    LocalMux I__5822 (
            .O(N__31831),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__5821 (
            .O(N__31828),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__5820 (
            .O(N__31823),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    CascadeMux I__5819 (
            .O(N__31820),
            .I(N__31816));
    CascadeMux I__5818 (
            .O(N__31819),
            .I(N__31813));
    InMux I__5817 (
            .O(N__31816),
            .I(N__31810));
    InMux I__5816 (
            .O(N__31813),
            .I(N__31807));
    LocalMux I__5815 (
            .O(N__31810),
            .I(N__31801));
    LocalMux I__5814 (
            .O(N__31807),
            .I(N__31801));
    InMux I__5813 (
            .O(N__31806),
            .I(N__31798));
    Span12Mux_s11_v I__5812 (
            .O(N__31801),
            .I(N__31795));
    LocalMux I__5811 (
            .O(N__31798),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv12 I__5810 (
            .O(N__31795),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__5809 (
            .O(N__31790),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    CascadeMux I__5808 (
            .O(N__31787),
            .I(N__31783));
    CascadeMux I__5807 (
            .O(N__31786),
            .I(N__31780));
    InMux I__5806 (
            .O(N__31783),
            .I(N__31774));
    InMux I__5805 (
            .O(N__31780),
            .I(N__31774));
    InMux I__5804 (
            .O(N__31779),
            .I(N__31771));
    LocalMux I__5803 (
            .O(N__31774),
            .I(N__31768));
    LocalMux I__5802 (
            .O(N__31771),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__5801 (
            .O(N__31768),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__5800 (
            .O(N__31763),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__5799 (
            .O(N__31760),
            .I(N__31754));
    InMux I__5798 (
            .O(N__31759),
            .I(N__31754));
    LocalMux I__5797 (
            .O(N__31754),
            .I(N__31750));
    InMux I__5796 (
            .O(N__31753),
            .I(N__31747));
    Span4Mux_v I__5795 (
            .O(N__31750),
            .I(N__31744));
    LocalMux I__5794 (
            .O(N__31747),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__5793 (
            .O(N__31744),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__5792 (
            .O(N__31739),
            .I(bfn_12_13_0_));
    CascadeMux I__5791 (
            .O(N__31736),
            .I(N__31733));
    InMux I__5790 (
            .O(N__31733),
            .I(N__31726));
    InMux I__5789 (
            .O(N__31732),
            .I(N__31726));
    InMux I__5788 (
            .O(N__31731),
            .I(N__31723));
    LocalMux I__5787 (
            .O(N__31726),
            .I(N__31720));
    LocalMux I__5786 (
            .O(N__31723),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv12 I__5785 (
            .O(N__31720),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__5784 (
            .O(N__31715),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__5783 (
            .O(N__31712),
            .I(N__31705));
    InMux I__5782 (
            .O(N__31711),
            .I(N__31705));
    InMux I__5781 (
            .O(N__31710),
            .I(N__31702));
    LocalMux I__5780 (
            .O(N__31705),
            .I(N__31699));
    LocalMux I__5779 (
            .O(N__31702),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__5778 (
            .O(N__31699),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__5777 (
            .O(N__31694),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    CascadeMux I__5776 (
            .O(N__31691),
            .I(N__31688));
    InMux I__5775 (
            .O(N__31688),
            .I(N__31681));
    InMux I__5774 (
            .O(N__31687),
            .I(N__31681));
    InMux I__5773 (
            .O(N__31686),
            .I(N__31678));
    LocalMux I__5772 (
            .O(N__31681),
            .I(N__31675));
    LocalMux I__5771 (
            .O(N__31678),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__5770 (
            .O(N__31675),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__5769 (
            .O(N__31670),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__5768 (
            .O(N__31667),
            .I(N__31664));
    LocalMux I__5767 (
            .O(N__31664),
            .I(N__31660));
    InMux I__5766 (
            .O(N__31663),
            .I(N__31657));
    Span4Mux_h I__5765 (
            .O(N__31660),
            .I(N__31654));
    LocalMux I__5764 (
            .O(N__31657),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__5763 (
            .O(N__31654),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__5762 (
            .O(N__31649),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__5761 (
            .O(N__31646),
            .I(N__31643));
    LocalMux I__5760 (
            .O(N__31643),
            .I(N__31639));
    InMux I__5759 (
            .O(N__31642),
            .I(N__31636));
    Span4Mux_h I__5758 (
            .O(N__31639),
            .I(N__31633));
    LocalMux I__5757 (
            .O(N__31636),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__5756 (
            .O(N__31633),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__5755 (
            .O(N__31628),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__5754 (
            .O(N__31625),
            .I(N__31622));
    LocalMux I__5753 (
            .O(N__31622),
            .I(N__31618));
    InMux I__5752 (
            .O(N__31621),
            .I(N__31615));
    Span4Mux_h I__5751 (
            .O(N__31618),
            .I(N__31612));
    LocalMux I__5750 (
            .O(N__31615),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__5749 (
            .O(N__31612),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__5748 (
            .O(N__31607),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__5747 (
            .O(N__31604),
            .I(N__31601));
    LocalMux I__5746 (
            .O(N__31601),
            .I(N__31597));
    InMux I__5745 (
            .O(N__31600),
            .I(N__31594));
    Span4Mux_h I__5744 (
            .O(N__31597),
            .I(N__31591));
    LocalMux I__5743 (
            .O(N__31594),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__5742 (
            .O(N__31591),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__5741 (
            .O(N__31586),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    CascadeMux I__5740 (
            .O(N__31583),
            .I(N__31580));
    InMux I__5739 (
            .O(N__31580),
            .I(N__31574));
    InMux I__5738 (
            .O(N__31579),
            .I(N__31574));
    LocalMux I__5737 (
            .O(N__31574),
            .I(N__31570));
    InMux I__5736 (
            .O(N__31573),
            .I(N__31567));
    Span4Mux_v I__5735 (
            .O(N__31570),
            .I(N__31564));
    LocalMux I__5734 (
            .O(N__31567),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__5733 (
            .O(N__31564),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__5732 (
            .O(N__31559),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__5731 (
            .O(N__31556),
            .I(N__31549));
    InMux I__5730 (
            .O(N__31555),
            .I(N__31549));
    InMux I__5729 (
            .O(N__31554),
            .I(N__31546));
    LocalMux I__5728 (
            .O(N__31549),
            .I(N__31543));
    LocalMux I__5727 (
            .O(N__31546),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__5726 (
            .O(N__31543),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__5725 (
            .O(N__31538),
            .I(bfn_12_12_0_));
    InMux I__5724 (
            .O(N__31535),
            .I(N__31529));
    InMux I__5723 (
            .O(N__31534),
            .I(N__31529));
    LocalMux I__5722 (
            .O(N__31529),
            .I(N__31526));
    Span4Mux_h I__5721 (
            .O(N__31526),
            .I(N__31522));
    InMux I__5720 (
            .O(N__31525),
            .I(N__31519));
    Span4Mux_v I__5719 (
            .O(N__31522),
            .I(N__31516));
    LocalMux I__5718 (
            .O(N__31519),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__5717 (
            .O(N__31516),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__5716 (
            .O(N__31511),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    CascadeMux I__5715 (
            .O(N__31508),
            .I(N__31504));
    InMux I__5714 (
            .O(N__31507),
            .I(N__31499));
    InMux I__5713 (
            .O(N__31504),
            .I(N__31499));
    LocalMux I__5712 (
            .O(N__31499),
            .I(N__31496));
    Span4Mux_v I__5711 (
            .O(N__31496),
            .I(N__31492));
    InMux I__5710 (
            .O(N__31495),
            .I(N__31489));
    Span4Mux_v I__5709 (
            .O(N__31492),
            .I(N__31486));
    LocalMux I__5708 (
            .O(N__31489),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__5707 (
            .O(N__31486),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__5706 (
            .O(N__31481),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__5705 (
            .O(N__31478),
            .I(N__31475));
    LocalMux I__5704 (
            .O(N__31475),
            .I(N__31471));
    InMux I__5703 (
            .O(N__31474),
            .I(N__31468));
    Span4Mux_h I__5702 (
            .O(N__31471),
            .I(N__31465));
    LocalMux I__5701 (
            .O(N__31468),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__5700 (
            .O(N__31465),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__5699 (
            .O(N__31460),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__5698 (
            .O(N__31457),
            .I(N__31454));
    LocalMux I__5697 (
            .O(N__31454),
            .I(N__31450));
    InMux I__5696 (
            .O(N__31453),
            .I(N__31447));
    Span4Mux_v I__5695 (
            .O(N__31450),
            .I(N__31444));
    LocalMux I__5694 (
            .O(N__31447),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__5693 (
            .O(N__31444),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__5692 (
            .O(N__31439),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__5691 (
            .O(N__31436),
            .I(N__31433));
    LocalMux I__5690 (
            .O(N__31433),
            .I(N__31429));
    InMux I__5689 (
            .O(N__31432),
            .I(N__31426));
    Span4Mux_v I__5688 (
            .O(N__31429),
            .I(N__31423));
    LocalMux I__5687 (
            .O(N__31426),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__5686 (
            .O(N__31423),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__5685 (
            .O(N__31418),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__5684 (
            .O(N__31415),
            .I(N__31412));
    LocalMux I__5683 (
            .O(N__31412),
            .I(N__31408));
    InMux I__5682 (
            .O(N__31411),
            .I(N__31405));
    Span4Mux_h I__5681 (
            .O(N__31408),
            .I(N__31402));
    LocalMux I__5680 (
            .O(N__31405),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__5679 (
            .O(N__31402),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__5678 (
            .O(N__31397),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__5677 (
            .O(N__31394),
            .I(N__31391));
    LocalMux I__5676 (
            .O(N__31391),
            .I(N__31387));
    InMux I__5675 (
            .O(N__31390),
            .I(N__31384));
    Span4Mux_h I__5674 (
            .O(N__31387),
            .I(N__31381));
    LocalMux I__5673 (
            .O(N__31384),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__5672 (
            .O(N__31381),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__5671 (
            .O(N__31376),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__5670 (
            .O(N__31373),
            .I(N__31370));
    LocalMux I__5669 (
            .O(N__31370),
            .I(N__31366));
    InMux I__5668 (
            .O(N__31369),
            .I(N__31363));
    Span4Mux_v I__5667 (
            .O(N__31366),
            .I(N__31360));
    LocalMux I__5666 (
            .O(N__31363),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__5665 (
            .O(N__31360),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__5664 (
            .O(N__31355),
            .I(bfn_12_11_0_));
    InMux I__5663 (
            .O(N__31352),
            .I(N__31349));
    LocalMux I__5662 (
            .O(N__31349),
            .I(N__31345));
    InMux I__5661 (
            .O(N__31348),
            .I(N__31342));
    Span4Mux_v I__5660 (
            .O(N__31345),
            .I(N__31339));
    LocalMux I__5659 (
            .O(N__31342),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__5658 (
            .O(N__31339),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__5657 (
            .O(N__31334),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__5656 (
            .O(N__31331),
            .I(N__31328));
    LocalMux I__5655 (
            .O(N__31328),
            .I(N__31324));
    InMux I__5654 (
            .O(N__31327),
            .I(N__31321));
    Span4Mux_h I__5653 (
            .O(N__31324),
            .I(N__31318));
    LocalMux I__5652 (
            .O(N__31321),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__5651 (
            .O(N__31318),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__5650 (
            .O(N__31313),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__5649 (
            .O(N__31310),
            .I(N__31306));
    InMux I__5648 (
            .O(N__31309),
            .I(N__31302));
    LocalMux I__5647 (
            .O(N__31306),
            .I(N__31299));
    InMux I__5646 (
            .O(N__31305),
            .I(N__31296));
    LocalMux I__5645 (
            .O(N__31302),
            .I(N__31289));
    Span12Mux_v I__5644 (
            .O(N__31299),
            .I(N__31289));
    LocalMux I__5643 (
            .O(N__31296),
            .I(N__31289));
    Odrv12 I__5642 (
            .O(N__31289),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    CascadeMux I__5641 (
            .O(N__31286),
            .I(N__31282));
    CascadeMux I__5640 (
            .O(N__31285),
            .I(N__31279));
    InMux I__5639 (
            .O(N__31282),
            .I(N__31276));
    InMux I__5638 (
            .O(N__31279),
            .I(N__31273));
    LocalMux I__5637 (
            .O(N__31276),
            .I(N__31270));
    LocalMux I__5636 (
            .O(N__31273),
            .I(N__31267));
    Span4Mux_v I__5635 (
            .O(N__31270),
            .I(N__31264));
    Span4Mux_h I__5634 (
            .O(N__31267),
            .I(N__31261));
    Odrv4 I__5633 (
            .O(N__31264),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    Odrv4 I__5632 (
            .O(N__31261),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    CascadeMux I__5631 (
            .O(N__31256),
            .I(N__31253));
    InMux I__5630 (
            .O(N__31253),
            .I(N__31250));
    LocalMux I__5629 (
            .O(N__31250),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    InMux I__5628 (
            .O(N__31247),
            .I(N__31244));
    LocalMux I__5627 (
            .O(N__31244),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    InMux I__5626 (
            .O(N__31241),
            .I(N__31238));
    LocalMux I__5625 (
            .O(N__31238),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__5624 (
            .O(N__31235),
            .I(N__31231));
    CascadeMux I__5623 (
            .O(N__31234),
            .I(N__31228));
    LocalMux I__5622 (
            .O(N__31231),
            .I(N__31225));
    InMux I__5621 (
            .O(N__31228),
            .I(N__31222));
    Span4Mux_v I__5620 (
            .O(N__31225),
            .I(N__31219));
    LocalMux I__5619 (
            .O(N__31222),
            .I(N__31214));
    Span4Mux_h I__5618 (
            .O(N__31219),
            .I(N__31211));
    InMux I__5617 (
            .O(N__31218),
            .I(N__31208));
    InMux I__5616 (
            .O(N__31217),
            .I(N__31205));
    Odrv12 I__5615 (
            .O(N__31214),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv4 I__5614 (
            .O(N__31211),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__5613 (
            .O(N__31208),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__5612 (
            .O(N__31205),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__5611 (
            .O(N__31196),
            .I(N__31193));
    LocalMux I__5610 (
            .O(N__31193),
            .I(N__31190));
    Span4Mux_v I__5609 (
            .O(N__31190),
            .I(N__31186));
    InMux I__5608 (
            .O(N__31189),
            .I(N__31183));
    Odrv4 I__5607 (
            .O(N__31186),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__5606 (
            .O(N__31183),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    InMux I__5605 (
            .O(N__31178),
            .I(N__31175));
    LocalMux I__5604 (
            .O(N__31175),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__5603 (
            .O(N__31172),
            .I(N__31168));
    InMux I__5602 (
            .O(N__31171),
            .I(N__31164));
    LocalMux I__5601 (
            .O(N__31168),
            .I(N__31161));
    CascadeMux I__5600 (
            .O(N__31167),
            .I(N__31158));
    LocalMux I__5599 (
            .O(N__31164),
            .I(N__31155));
    Span4Mux_v I__5598 (
            .O(N__31161),
            .I(N__31152));
    InMux I__5597 (
            .O(N__31158),
            .I(N__31149));
    Span12Mux_h I__5596 (
            .O(N__31155),
            .I(N__31146));
    Span4Mux_h I__5595 (
            .O(N__31152),
            .I(N__31143));
    LocalMux I__5594 (
            .O(N__31149),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__5593 (
            .O(N__31146),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__5592 (
            .O(N__31143),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__5591 (
            .O(N__31136),
            .I(N__31133));
    InMux I__5590 (
            .O(N__31133),
            .I(N__31130));
    LocalMux I__5589 (
            .O(N__31130),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    InMux I__5588 (
            .O(N__31127),
            .I(N__31124));
    LocalMux I__5587 (
            .O(N__31124),
            .I(N__31120));
    InMux I__5586 (
            .O(N__31123),
            .I(N__31117));
    Span4Mux_v I__5585 (
            .O(N__31120),
            .I(N__31114));
    LocalMux I__5584 (
            .O(N__31117),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__5583 (
            .O(N__31114),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__5582 (
            .O(N__31109),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__5581 (
            .O(N__31106),
            .I(N__31103));
    LocalMux I__5580 (
            .O(N__31103),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ));
    InMux I__5579 (
            .O(N__31100),
            .I(N__31096));
    CascadeMux I__5578 (
            .O(N__31099),
            .I(N__31093));
    LocalMux I__5577 (
            .O(N__31096),
            .I(N__31090));
    InMux I__5576 (
            .O(N__31093),
            .I(N__31087));
    Span4Mux_h I__5575 (
            .O(N__31090),
            .I(N__31084));
    LocalMux I__5574 (
            .O(N__31087),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__5573 (
            .O(N__31084),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__5572 (
            .O(N__31079),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__5571 (
            .O(N__31076),
            .I(N__31073));
    LocalMux I__5570 (
            .O(N__31073),
            .I(N__31068));
    InMux I__5569 (
            .O(N__31072),
            .I(N__31065));
    InMux I__5568 (
            .O(N__31071),
            .I(N__31062));
    Span4Mux_v I__5567 (
            .O(N__31068),
            .I(N__31059));
    LocalMux I__5566 (
            .O(N__31065),
            .I(N__31056));
    LocalMux I__5565 (
            .O(N__31062),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__5564 (
            .O(N__31059),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__5563 (
            .O(N__31056),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    CascadeMux I__5562 (
            .O(N__31049),
            .I(N__31043));
    InMux I__5561 (
            .O(N__31048),
            .I(N__31036));
    InMux I__5560 (
            .O(N__31047),
            .I(N__31036));
    InMux I__5559 (
            .O(N__31046),
            .I(N__31036));
    InMux I__5558 (
            .O(N__31043),
            .I(N__31033));
    LocalMux I__5557 (
            .O(N__31036),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5556 (
            .O(N__31033),
            .I(\phase_controller_inst1.hc_time_passed ));
    CascadeMux I__5555 (
            .O(N__31028),
            .I(N__31024));
    InMux I__5554 (
            .O(N__31027),
            .I(N__31015));
    InMux I__5553 (
            .O(N__31024),
            .I(N__31015));
    InMux I__5552 (
            .O(N__31023),
            .I(N__31015));
    InMux I__5551 (
            .O(N__31022),
            .I(N__31012));
    LocalMux I__5550 (
            .O(N__31015),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__5549 (
            .O(N__31012),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    IoInMux I__5548 (
            .O(N__31007),
            .I(N__31004));
    LocalMux I__5547 (
            .O(N__31004),
            .I(N__31001));
    IoSpan4Mux I__5546 (
            .O(N__31001),
            .I(N__30998));
    Span4Mux_s0_v I__5545 (
            .O(N__30998),
            .I(N__30995));
    Sp12to4 I__5544 (
            .O(N__30995),
            .I(N__30992));
    Span12Mux_v I__5543 (
            .O(N__30992),
            .I(N__30989));
    Span12Mux_v I__5542 (
            .O(N__30989),
            .I(N__30985));
    InMux I__5541 (
            .O(N__30988),
            .I(N__30982));
    Odrv12 I__5540 (
            .O(N__30985),
            .I(test22_c));
    LocalMux I__5539 (
            .O(N__30982),
            .I(test22_c));
    InMux I__5538 (
            .O(N__30977),
            .I(N__30974));
    LocalMux I__5537 (
            .O(N__30974),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    InMux I__5536 (
            .O(N__30971),
            .I(N__30968));
    LocalMux I__5535 (
            .O(N__30968),
            .I(N__30964));
    InMux I__5534 (
            .O(N__30967),
            .I(N__30961));
    Span4Mux_s3_h I__5533 (
            .O(N__30964),
            .I(N__30958));
    LocalMux I__5532 (
            .O(N__30961),
            .I(N__30955));
    Span4Mux_v I__5531 (
            .O(N__30958),
            .I(N__30952));
    Span12Mux_s8_h I__5530 (
            .O(N__30955),
            .I(N__30947));
    Sp12to4 I__5529 (
            .O(N__30952),
            .I(N__30947));
    Odrv12 I__5528 (
            .O(N__30947),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__5527 (
            .O(N__30944),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__5526 (
            .O(N__30941),
            .I(N__30938));
    LocalMux I__5525 (
            .O(N__30938),
            .I(N__30935));
    Span4Mux_v I__5524 (
            .O(N__30935),
            .I(N__30932));
    Span4Mux_h I__5523 (
            .O(N__30932),
            .I(N__30929));
    Span4Mux_h I__5522 (
            .O(N__30929),
            .I(N__30925));
    InMux I__5521 (
            .O(N__30928),
            .I(N__30922));
    Span4Mux_h I__5520 (
            .O(N__30925),
            .I(N__30919));
    LocalMux I__5519 (
            .O(N__30922),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    Odrv4 I__5518 (
            .O(N__30919),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__5517 (
            .O(N__30914),
            .I(bfn_11_22_0_));
    InMux I__5516 (
            .O(N__30911),
            .I(N__30908));
    LocalMux I__5515 (
            .O(N__30908),
            .I(N__30905));
    Span4Mux_v I__5514 (
            .O(N__30905),
            .I(N__30902));
    Span4Mux_h I__5513 (
            .O(N__30902),
            .I(N__30898));
    InMux I__5512 (
            .O(N__30901),
            .I(N__30895));
    Span4Mux_h I__5511 (
            .O(N__30898),
            .I(N__30892));
    LocalMux I__5510 (
            .O(N__30895),
            .I(N__30887));
    Span4Mux_h I__5509 (
            .O(N__30892),
            .I(N__30887));
    Odrv4 I__5508 (
            .O(N__30887),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__5507 (
            .O(N__30884),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__5506 (
            .O(N__30881),
            .I(N__30878));
    LocalMux I__5505 (
            .O(N__30878),
            .I(N__30875));
    Span4Mux_s1_h I__5504 (
            .O(N__30875),
            .I(N__30872));
    Span4Mux_h I__5503 (
            .O(N__30872),
            .I(N__30868));
    InMux I__5502 (
            .O(N__30871),
            .I(N__30865));
    Span4Mux_h I__5501 (
            .O(N__30868),
            .I(N__30862));
    LocalMux I__5500 (
            .O(N__30865),
            .I(N__30859));
    Span4Mux_h I__5499 (
            .O(N__30862),
            .I(N__30856));
    Odrv4 I__5498 (
            .O(N__30859),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv4 I__5497 (
            .O(N__30856),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__5496 (
            .O(N__30851),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__5495 (
            .O(N__30848),
            .I(N__30845));
    LocalMux I__5494 (
            .O(N__30845),
            .I(N__30841));
    InMux I__5493 (
            .O(N__30844),
            .I(N__30838));
    Span12Mux_s2_h I__5492 (
            .O(N__30841),
            .I(N__30835));
    LocalMux I__5491 (
            .O(N__30838),
            .I(N__30832));
    Span12Mux_h I__5490 (
            .O(N__30835),
            .I(N__30829));
    Odrv4 I__5489 (
            .O(N__30832),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    Odrv12 I__5488 (
            .O(N__30829),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    InMux I__5487 (
            .O(N__30824),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ));
    InMux I__5486 (
            .O(N__30821),
            .I(N__30818));
    LocalMux I__5485 (
            .O(N__30818),
            .I(N__30815));
    Span4Mux_s1_h I__5484 (
            .O(N__30815),
            .I(N__30812));
    Span4Mux_h I__5483 (
            .O(N__30812),
            .I(N__30809));
    Span4Mux_h I__5482 (
            .O(N__30809),
            .I(N__30805));
    InMux I__5481 (
            .O(N__30808),
            .I(N__30802));
    Span4Mux_h I__5480 (
            .O(N__30805),
            .I(N__30799));
    LocalMux I__5479 (
            .O(N__30802),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    Odrv4 I__5478 (
            .O(N__30799),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    InMux I__5477 (
            .O(N__30794),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ));
    InMux I__5476 (
            .O(N__30791),
            .I(N__30788));
    LocalMux I__5475 (
            .O(N__30788),
            .I(N__30785));
    Span4Mux_s3_h I__5474 (
            .O(N__30785),
            .I(N__30781));
    InMux I__5473 (
            .O(N__30784),
            .I(N__30778));
    Sp12to4 I__5472 (
            .O(N__30781),
            .I(N__30775));
    LocalMux I__5471 (
            .O(N__30778),
            .I(N__30770));
    Span12Mux_s8_v I__5470 (
            .O(N__30775),
            .I(N__30770));
    Odrv12 I__5469 (
            .O(N__30770),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    InMux I__5468 (
            .O(N__30767),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ));
    InMux I__5467 (
            .O(N__30764),
            .I(N__30761));
    LocalMux I__5466 (
            .O(N__30761),
            .I(N__30758));
    Span12Mux_s8_v I__5465 (
            .O(N__30758),
            .I(N__30754));
    InMux I__5464 (
            .O(N__30757),
            .I(N__30751));
    Span12Mux_h I__5463 (
            .O(N__30754),
            .I(N__30748));
    LocalMux I__5462 (
            .O(N__30751),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    Odrv12 I__5461 (
            .O(N__30748),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    InMux I__5460 (
            .O(N__30743),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ));
    InMux I__5459 (
            .O(N__30740),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ));
    InMux I__5458 (
            .O(N__30737),
            .I(N__30734));
    LocalMux I__5457 (
            .O(N__30734),
            .I(N__30731));
    Odrv4 I__5456 (
            .O(N__30731),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_31 ));
    InMux I__5455 (
            .O(N__30728),
            .I(N__30725));
    LocalMux I__5454 (
            .O(N__30725),
            .I(N__30722));
    Span4Mux_v I__5453 (
            .O(N__30722),
            .I(N__30718));
    InMux I__5452 (
            .O(N__30721),
            .I(N__30715));
    Sp12to4 I__5451 (
            .O(N__30718),
            .I(N__30712));
    LocalMux I__5450 (
            .O(N__30715),
            .I(N__30709));
    Span12Mux_h I__5449 (
            .O(N__30712),
            .I(N__30706));
    Odrv4 I__5448 (
            .O(N__30709),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    Odrv12 I__5447 (
            .O(N__30706),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__5446 (
            .O(N__30701),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__5445 (
            .O(N__30698),
            .I(N__30695));
    LocalMux I__5444 (
            .O(N__30695),
            .I(N__30692));
    Span4Mux_s2_h I__5443 (
            .O(N__30692),
            .I(N__30688));
    InMux I__5442 (
            .O(N__30691),
            .I(N__30685));
    Span4Mux_h I__5441 (
            .O(N__30688),
            .I(N__30682));
    LocalMux I__5440 (
            .O(N__30685),
            .I(N__30679));
    Span4Mux_h I__5439 (
            .O(N__30682),
            .I(N__30676));
    Span4Mux_v I__5438 (
            .O(N__30679),
            .I(N__30673));
    Span4Mux_v I__5437 (
            .O(N__30676),
            .I(N__30670));
    Odrv4 I__5436 (
            .O(N__30673),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv4 I__5435 (
            .O(N__30670),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__5434 (
            .O(N__30665),
            .I(bfn_11_21_0_));
    InMux I__5433 (
            .O(N__30662),
            .I(N__30659));
    LocalMux I__5432 (
            .O(N__30659),
            .I(N__30656));
    Span4Mux_v I__5431 (
            .O(N__30656),
            .I(N__30652));
    InMux I__5430 (
            .O(N__30655),
            .I(N__30649));
    Sp12to4 I__5429 (
            .O(N__30652),
            .I(N__30646));
    LocalMux I__5428 (
            .O(N__30649),
            .I(N__30643));
    Span12Mux_h I__5427 (
            .O(N__30646),
            .I(N__30640));
    Odrv12 I__5426 (
            .O(N__30643),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    Odrv12 I__5425 (
            .O(N__30640),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__5424 (
            .O(N__30635),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__5423 (
            .O(N__30632),
            .I(N__30629));
    LocalMux I__5422 (
            .O(N__30629),
            .I(N__30626));
    Span4Mux_s2_h I__5421 (
            .O(N__30626),
            .I(N__30623));
    Span4Mux_h I__5420 (
            .O(N__30623),
            .I(N__30619));
    InMux I__5419 (
            .O(N__30622),
            .I(N__30616));
    Span4Mux_h I__5418 (
            .O(N__30619),
            .I(N__30613));
    LocalMux I__5417 (
            .O(N__30616),
            .I(N__30610));
    Span4Mux_v I__5416 (
            .O(N__30613),
            .I(N__30607));
    Odrv4 I__5415 (
            .O(N__30610),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    Odrv4 I__5414 (
            .O(N__30607),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__5413 (
            .O(N__30602),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__5412 (
            .O(N__30599),
            .I(N__30596));
    LocalMux I__5411 (
            .O(N__30596),
            .I(N__30593));
    Span4Mux_v I__5410 (
            .O(N__30593),
            .I(N__30589));
    InMux I__5409 (
            .O(N__30592),
            .I(N__30586));
    Sp12to4 I__5408 (
            .O(N__30589),
            .I(N__30583));
    LocalMux I__5407 (
            .O(N__30586),
            .I(N__30580));
    Span12Mux_h I__5406 (
            .O(N__30583),
            .I(N__30577));
    Odrv12 I__5405 (
            .O(N__30580),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    Odrv12 I__5404 (
            .O(N__30577),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    InMux I__5403 (
            .O(N__30572),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__5402 (
            .O(N__30569),
            .I(N__30566));
    LocalMux I__5401 (
            .O(N__30566),
            .I(N__30562));
    InMux I__5400 (
            .O(N__30565),
            .I(N__30559));
    Span12Mux_s2_h I__5399 (
            .O(N__30562),
            .I(N__30556));
    LocalMux I__5398 (
            .O(N__30559),
            .I(N__30553));
    Span12Mux_h I__5397 (
            .O(N__30556),
            .I(N__30550));
    Odrv4 I__5396 (
            .O(N__30553),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    Odrv12 I__5395 (
            .O(N__30550),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    InMux I__5394 (
            .O(N__30545),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__5393 (
            .O(N__30542),
            .I(N__30539));
    LocalMux I__5392 (
            .O(N__30539),
            .I(N__30536));
    Span4Mux_s1_h I__5391 (
            .O(N__30536),
            .I(N__30532));
    InMux I__5390 (
            .O(N__30535),
            .I(N__30529));
    Span4Mux_v I__5389 (
            .O(N__30532),
            .I(N__30526));
    LocalMux I__5388 (
            .O(N__30529),
            .I(N__30523));
    Sp12to4 I__5387 (
            .O(N__30526),
            .I(N__30520));
    Odrv4 I__5386 (
            .O(N__30523),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    Odrv12 I__5385 (
            .O(N__30520),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__5384 (
            .O(N__30515),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__5383 (
            .O(N__30512),
            .I(N__30509));
    LocalMux I__5382 (
            .O(N__30509),
            .I(N__30505));
    InMux I__5381 (
            .O(N__30508),
            .I(N__30502));
    Span12Mux_s9_v I__5380 (
            .O(N__30505),
            .I(N__30499));
    LocalMux I__5379 (
            .O(N__30502),
            .I(N__30494));
    Span12Mux_h I__5378 (
            .O(N__30499),
            .I(N__30494));
    Odrv12 I__5377 (
            .O(N__30494),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    InMux I__5376 (
            .O(N__30491),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    InMux I__5375 (
            .O(N__30488),
            .I(N__30485));
    LocalMux I__5374 (
            .O(N__30485),
            .I(N__30482));
    Span4Mux_s3_h I__5373 (
            .O(N__30482),
            .I(N__30478));
    InMux I__5372 (
            .O(N__30481),
            .I(N__30475));
    Span4Mux_h I__5371 (
            .O(N__30478),
            .I(N__30472));
    LocalMux I__5370 (
            .O(N__30475),
            .I(N__30469));
    Span4Mux_h I__5369 (
            .O(N__30472),
            .I(N__30466));
    Span12Mux_s9_h I__5368 (
            .O(N__30469),
            .I(N__30463));
    Span4Mux_v I__5367 (
            .O(N__30466),
            .I(N__30460));
    Odrv12 I__5366 (
            .O(N__30463),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__5365 (
            .O(N__30460),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__5364 (
            .O(N__30455),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__5363 (
            .O(N__30452),
            .I(N__30449));
    LocalMux I__5362 (
            .O(N__30449),
            .I(N__30445));
    InMux I__5361 (
            .O(N__30448),
            .I(N__30442));
    Span4Mux_h I__5360 (
            .O(N__30445),
            .I(N__30439));
    LocalMux I__5359 (
            .O(N__30442),
            .I(N__30436));
    Span4Mux_h I__5358 (
            .O(N__30439),
            .I(N__30433));
    Span12Mux_v I__5357 (
            .O(N__30436),
            .I(N__30430));
    Odrv4 I__5356 (
            .O(N__30433),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv12 I__5355 (
            .O(N__30430),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__5354 (
            .O(N__30425),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__5353 (
            .O(N__30422),
            .I(N__30418));
    InMux I__5352 (
            .O(N__30421),
            .I(N__30415));
    LocalMux I__5351 (
            .O(N__30418),
            .I(N__30412));
    LocalMux I__5350 (
            .O(N__30415),
            .I(N__30409));
    Span4Mux_h I__5349 (
            .O(N__30412),
            .I(N__30406));
    Span4Mux_v I__5348 (
            .O(N__30409),
            .I(N__30401));
    Span4Mux_v I__5347 (
            .O(N__30406),
            .I(N__30401));
    Sp12to4 I__5346 (
            .O(N__30401),
            .I(N__30398));
    Span12Mux_s11_h I__5345 (
            .O(N__30398),
            .I(N__30395));
    Odrv12 I__5344 (
            .O(N__30395),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__5343 (
            .O(N__30392),
            .I(bfn_11_20_0_));
    InMux I__5342 (
            .O(N__30389),
            .I(N__30386));
    LocalMux I__5341 (
            .O(N__30386),
            .I(N__30383));
    Span4Mux_v I__5340 (
            .O(N__30383),
            .I(N__30380));
    Sp12to4 I__5339 (
            .O(N__30380),
            .I(N__30376));
    InMux I__5338 (
            .O(N__30379),
            .I(N__30373));
    Span12Mux_s6_h I__5337 (
            .O(N__30376),
            .I(N__30370));
    LocalMux I__5336 (
            .O(N__30373),
            .I(N__30365));
    Span12Mux_v I__5335 (
            .O(N__30370),
            .I(N__30365));
    Odrv12 I__5334 (
            .O(N__30365),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__5333 (
            .O(N__30362),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__5332 (
            .O(N__30359),
            .I(N__30356));
    LocalMux I__5331 (
            .O(N__30356),
            .I(N__30353));
    Span4Mux_v I__5330 (
            .O(N__30353),
            .I(N__30349));
    InMux I__5329 (
            .O(N__30352),
            .I(N__30346));
    Sp12to4 I__5328 (
            .O(N__30349),
            .I(N__30343));
    LocalMux I__5327 (
            .O(N__30346),
            .I(N__30340));
    Span12Mux_s11_h I__5326 (
            .O(N__30343),
            .I(N__30337));
    Odrv12 I__5325 (
            .O(N__30340),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv12 I__5324 (
            .O(N__30337),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__5323 (
            .O(N__30332),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__5322 (
            .O(N__30329),
            .I(N__30326));
    LocalMux I__5321 (
            .O(N__30326),
            .I(N__30323));
    Span4Mux_v I__5320 (
            .O(N__30323),
            .I(N__30319));
    InMux I__5319 (
            .O(N__30322),
            .I(N__30316));
    Sp12to4 I__5318 (
            .O(N__30319),
            .I(N__30313));
    LocalMux I__5317 (
            .O(N__30316),
            .I(N__30310));
    Span12Mux_s11_h I__5316 (
            .O(N__30313),
            .I(N__30307));
    Odrv12 I__5315 (
            .O(N__30310),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv12 I__5314 (
            .O(N__30307),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__5313 (
            .O(N__30302),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__5312 (
            .O(N__30299),
            .I(N__30295));
    InMux I__5311 (
            .O(N__30298),
            .I(N__30292));
    LocalMux I__5310 (
            .O(N__30295),
            .I(N__30289));
    LocalMux I__5309 (
            .O(N__30292),
            .I(N__30286));
    Span12Mux_s11_h I__5308 (
            .O(N__30289),
            .I(N__30283));
    Odrv12 I__5307 (
            .O(N__30286),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv12 I__5306 (
            .O(N__30283),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__5305 (
            .O(N__30278),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__5304 (
            .O(N__30275),
            .I(N__30272));
    LocalMux I__5303 (
            .O(N__30272),
            .I(N__30269));
    Span4Mux_s3_h I__5302 (
            .O(N__30269),
            .I(N__30265));
    InMux I__5301 (
            .O(N__30268),
            .I(N__30262));
    Span4Mux_v I__5300 (
            .O(N__30265),
            .I(N__30259));
    LocalMux I__5299 (
            .O(N__30262),
            .I(N__30256));
    Span4Mux_h I__5298 (
            .O(N__30259),
            .I(N__30253));
    Span4Mux_h I__5297 (
            .O(N__30256),
            .I(N__30248));
    Span4Mux_h I__5296 (
            .O(N__30253),
            .I(N__30248));
    Odrv4 I__5295 (
            .O(N__30248),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__5294 (
            .O(N__30245),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__5293 (
            .O(N__30242),
            .I(N__30239));
    LocalMux I__5292 (
            .O(N__30239),
            .I(N__30236));
    Span4Mux_v I__5291 (
            .O(N__30236),
            .I(N__30232));
    InMux I__5290 (
            .O(N__30235),
            .I(N__30229));
    Sp12to4 I__5289 (
            .O(N__30232),
            .I(N__30226));
    LocalMux I__5288 (
            .O(N__30229),
            .I(N__30223));
    Span12Mux_s11_h I__5287 (
            .O(N__30226),
            .I(N__30220));
    Odrv12 I__5286 (
            .O(N__30223),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv12 I__5285 (
            .O(N__30220),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__5284 (
            .O(N__30215),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__5283 (
            .O(N__30212),
            .I(N__30209));
    LocalMux I__5282 (
            .O(N__30209),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__5281 (
            .O(N__30206),
            .I(N__30203));
    LocalMux I__5280 (
            .O(N__30203),
            .I(N__30200));
    Span4Mux_s3_h I__5279 (
            .O(N__30200),
            .I(N__30196));
    InMux I__5278 (
            .O(N__30199),
            .I(N__30193));
    Span4Mux_v I__5277 (
            .O(N__30196),
            .I(N__30190));
    LocalMux I__5276 (
            .O(N__30193),
            .I(N__30187));
    Span4Mux_h I__5275 (
            .O(N__30190),
            .I(N__30184));
    Span12Mux_s6_h I__5274 (
            .O(N__30187),
            .I(N__30181));
    Span4Mux_h I__5273 (
            .O(N__30184),
            .I(N__30178));
    Odrv12 I__5272 (
            .O(N__30181),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    Odrv4 I__5271 (
            .O(N__30178),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__5270 (
            .O(N__30173),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__5269 (
            .O(N__30170),
            .I(N__30167));
    LocalMux I__5268 (
            .O(N__30167),
            .I(N__30163));
    InMux I__5267 (
            .O(N__30166),
            .I(N__30160));
    Span4Mux_v I__5266 (
            .O(N__30163),
            .I(N__30157));
    LocalMux I__5265 (
            .O(N__30160),
            .I(N__30154));
    Sp12to4 I__5264 (
            .O(N__30157),
            .I(N__30151));
    Span12Mux_v I__5263 (
            .O(N__30154),
            .I(N__30148));
    Span12Mux_s11_h I__5262 (
            .O(N__30151),
            .I(N__30145));
    Odrv12 I__5261 (
            .O(N__30148),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv12 I__5260 (
            .O(N__30145),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__5259 (
            .O(N__30140),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__5258 (
            .O(N__30137),
            .I(N__30134));
    LocalMux I__5257 (
            .O(N__30134),
            .I(N__30130));
    InMux I__5256 (
            .O(N__30133),
            .I(N__30127));
    Span4Mux_h I__5255 (
            .O(N__30130),
            .I(N__30124));
    LocalMux I__5254 (
            .O(N__30127),
            .I(N__30121));
    Sp12to4 I__5253 (
            .O(N__30124),
            .I(N__30118));
    Span12Mux_s4_h I__5252 (
            .O(N__30121),
            .I(N__30113));
    Span12Mux_v I__5251 (
            .O(N__30118),
            .I(N__30113));
    Odrv12 I__5250 (
            .O(N__30113),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__5249 (
            .O(N__30110),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__5248 (
            .O(N__30107),
            .I(N__30103));
    InMux I__5247 (
            .O(N__30106),
            .I(N__30100));
    LocalMux I__5246 (
            .O(N__30103),
            .I(N__30097));
    LocalMux I__5245 (
            .O(N__30100),
            .I(N__30094));
    Span4Mux_v I__5244 (
            .O(N__30097),
            .I(N__30091));
    Span4Mux_h I__5243 (
            .O(N__30094),
            .I(N__30088));
    Sp12to4 I__5242 (
            .O(N__30091),
            .I(N__30085));
    Span4Mux_h I__5241 (
            .O(N__30088),
            .I(N__30082));
    Span12Mux_s11_h I__5240 (
            .O(N__30085),
            .I(N__30079));
    Odrv4 I__5239 (
            .O(N__30082),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv12 I__5238 (
            .O(N__30079),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__5237 (
            .O(N__30074),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__5236 (
            .O(N__30071),
            .I(N__30067));
    InMux I__5235 (
            .O(N__30070),
            .I(N__30064));
    LocalMux I__5234 (
            .O(N__30067),
            .I(N__30061));
    LocalMux I__5233 (
            .O(N__30064),
            .I(N__30058));
    Span4Mux_s2_h I__5232 (
            .O(N__30061),
            .I(N__30055));
    Span4Mux_v I__5231 (
            .O(N__30058),
            .I(N__30052));
    Sp12to4 I__5230 (
            .O(N__30055),
            .I(N__30049));
    Sp12to4 I__5229 (
            .O(N__30052),
            .I(N__30044));
    Span12Mux_v I__5228 (
            .O(N__30049),
            .I(N__30044));
    Odrv12 I__5227 (
            .O(N__30044),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__5226 (
            .O(N__30041),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    CascadeMux I__5225 (
            .O(N__30038),
            .I(N__30034));
    InMux I__5224 (
            .O(N__30037),
            .I(N__30028));
    InMux I__5223 (
            .O(N__30034),
            .I(N__30028));
    InMux I__5222 (
            .O(N__30033),
            .I(N__30025));
    LocalMux I__5221 (
            .O(N__30028),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__5220 (
            .O(N__30025),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__5219 (
            .O(N__30020),
            .I(N__30016));
    InMux I__5218 (
            .O(N__30019),
            .I(N__30013));
    LocalMux I__5217 (
            .O(N__30016),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__5216 (
            .O(N__30013),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__5215 (
            .O(N__30008),
            .I(N__30004));
    InMux I__5214 (
            .O(N__30007),
            .I(N__30001));
    LocalMux I__5213 (
            .O(N__30004),
            .I(N__29996));
    LocalMux I__5212 (
            .O(N__30001),
            .I(N__29996));
    Span4Mux_s3_v I__5211 (
            .O(N__29996),
            .I(N__29991));
    InMux I__5210 (
            .O(N__29995),
            .I(N__29988));
    InMux I__5209 (
            .O(N__29994),
            .I(N__29985));
    Span4Mux_h I__5208 (
            .O(N__29991),
            .I(N__29982));
    LocalMux I__5207 (
            .O(N__29988),
            .I(N__29979));
    LocalMux I__5206 (
            .O(N__29985),
            .I(N__29976));
    Sp12to4 I__5205 (
            .O(N__29982),
            .I(N__29973));
    Span4Mux_h I__5204 (
            .O(N__29979),
            .I(N__29970));
    Span4Mux_v I__5203 (
            .O(N__29976),
            .I(N__29967));
    Span12Mux_s11_v I__5202 (
            .O(N__29973),
            .I(N__29962));
    Sp12to4 I__5201 (
            .O(N__29970),
            .I(N__29962));
    Span4Mux_v I__5200 (
            .O(N__29967),
            .I(N__29959));
    Span12Mux_v I__5199 (
            .O(N__29962),
            .I(N__29956));
    Sp12to4 I__5198 (
            .O(N__29959),
            .I(N__29953));
    Span12Mux_h I__5197 (
            .O(N__29956),
            .I(N__29950));
    Span12Mux_h I__5196 (
            .O(N__29953),
            .I(N__29947));
    Odrv12 I__5195 (
            .O(N__29950),
            .I(start_stop_c));
    Odrv12 I__5194 (
            .O(N__29947),
            .I(start_stop_c));
    InMux I__5193 (
            .O(N__29942),
            .I(N__29939));
    LocalMux I__5192 (
            .O(N__29939),
            .I(N__29936));
    Span4Mux_v I__5191 (
            .O(N__29936),
            .I(N__29931));
    InMux I__5190 (
            .O(N__29935),
            .I(N__29928));
    InMux I__5189 (
            .O(N__29934),
            .I(N__29925));
    Sp12to4 I__5188 (
            .O(N__29931),
            .I(N__29918));
    LocalMux I__5187 (
            .O(N__29928),
            .I(N__29918));
    LocalMux I__5186 (
            .O(N__29925),
            .I(N__29918));
    Span12Mux_h I__5185 (
            .O(N__29918),
            .I(N__29915));
    Span12Mux_v I__5184 (
            .O(N__29915),
            .I(N__29912));
    Odrv12 I__5183 (
            .O(N__29912),
            .I(il_max_comp2_c));
    CascadeMux I__5182 (
            .O(N__29909),
            .I(phase_controller_inst1_N_54_cascade_));
    InMux I__5181 (
            .O(N__29906),
            .I(N__29903));
    LocalMux I__5180 (
            .O(N__29903),
            .I(N__29899));
    InMux I__5179 (
            .O(N__29902),
            .I(N__29896));
    Odrv4 I__5178 (
            .O(N__29899),
            .I(\phase_controller_inst2.N_54 ));
    LocalMux I__5177 (
            .O(N__29896),
            .I(\phase_controller_inst2.N_54 ));
    CascadeMux I__5176 (
            .O(N__29891),
            .I(N__29888));
    InMux I__5175 (
            .O(N__29888),
            .I(N__29884));
    InMux I__5174 (
            .O(N__29887),
            .I(N__29881));
    LocalMux I__5173 (
            .O(N__29884),
            .I(N__29875));
    LocalMux I__5172 (
            .O(N__29881),
            .I(N__29875));
    InMux I__5171 (
            .O(N__29880),
            .I(N__29871));
    Span12Mux_v I__5170 (
            .O(N__29875),
            .I(N__29868));
    InMux I__5169 (
            .O(N__29874),
            .I(N__29865));
    LocalMux I__5168 (
            .O(N__29871),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__5167 (
            .O(N__29868),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__5166 (
            .O(N__29865),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    CEMux I__5165 (
            .O(N__29858),
            .I(N__29853));
    CEMux I__5164 (
            .O(N__29857),
            .I(N__29849));
    CEMux I__5163 (
            .O(N__29856),
            .I(N__29846));
    LocalMux I__5162 (
            .O(N__29853),
            .I(N__29843));
    CEMux I__5161 (
            .O(N__29852),
            .I(N__29840));
    LocalMux I__5160 (
            .O(N__29849),
            .I(N__29837));
    LocalMux I__5159 (
            .O(N__29846),
            .I(N__29834));
    Span4Mux_v I__5158 (
            .O(N__29843),
            .I(N__29829));
    LocalMux I__5157 (
            .O(N__29840),
            .I(N__29829));
    Span4Mux_v I__5156 (
            .O(N__29837),
            .I(N__29826));
    Span4Mux_v I__5155 (
            .O(N__29834),
            .I(N__29823));
    Span4Mux_h I__5154 (
            .O(N__29829),
            .I(N__29820));
    Odrv4 I__5153 (
            .O(N__29826),
            .I(\delay_measurement_inst.delay_tr_timer.N_166_i ));
    Odrv4 I__5152 (
            .O(N__29823),
            .I(\delay_measurement_inst.delay_tr_timer.N_166_i ));
    Odrv4 I__5151 (
            .O(N__29820),
            .I(\delay_measurement_inst.delay_tr_timer.N_166_i ));
    CascadeMux I__5150 (
            .O(N__29813),
            .I(N__29809));
    InMux I__5149 (
            .O(N__29812),
            .I(N__29804));
    InMux I__5148 (
            .O(N__29809),
            .I(N__29799));
    InMux I__5147 (
            .O(N__29808),
            .I(N__29799));
    InMux I__5146 (
            .O(N__29807),
            .I(N__29796));
    LocalMux I__5145 (
            .O(N__29804),
            .I(N__29793));
    LocalMux I__5144 (
            .O(N__29799),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__5143 (
            .O(N__29796),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__5142 (
            .O(N__29793),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__5141 (
            .O(N__29786),
            .I(N__29780));
    InMux I__5140 (
            .O(N__29785),
            .I(N__29777));
    InMux I__5139 (
            .O(N__29784),
            .I(N__29772));
    InMux I__5138 (
            .O(N__29783),
            .I(N__29772));
    LocalMux I__5137 (
            .O(N__29780),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__5136 (
            .O(N__29777),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__5135 (
            .O(N__29772),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__5134 (
            .O(N__29765),
            .I(N__29753));
    InMux I__5133 (
            .O(N__29764),
            .I(N__29753));
    InMux I__5132 (
            .O(N__29763),
            .I(N__29753));
    InMux I__5131 (
            .O(N__29762),
            .I(N__29753));
    LocalMux I__5130 (
            .O(N__29753),
            .I(N__29728));
    InMux I__5129 (
            .O(N__29752),
            .I(N__29719));
    InMux I__5128 (
            .O(N__29751),
            .I(N__29719));
    InMux I__5127 (
            .O(N__29750),
            .I(N__29719));
    InMux I__5126 (
            .O(N__29749),
            .I(N__29719));
    InMux I__5125 (
            .O(N__29748),
            .I(N__29710));
    InMux I__5124 (
            .O(N__29747),
            .I(N__29710));
    InMux I__5123 (
            .O(N__29746),
            .I(N__29710));
    InMux I__5122 (
            .O(N__29745),
            .I(N__29710));
    InMux I__5121 (
            .O(N__29744),
            .I(N__29701));
    InMux I__5120 (
            .O(N__29743),
            .I(N__29701));
    InMux I__5119 (
            .O(N__29742),
            .I(N__29692));
    InMux I__5118 (
            .O(N__29741),
            .I(N__29692));
    InMux I__5117 (
            .O(N__29740),
            .I(N__29692));
    InMux I__5116 (
            .O(N__29739),
            .I(N__29692));
    InMux I__5115 (
            .O(N__29738),
            .I(N__29683));
    InMux I__5114 (
            .O(N__29737),
            .I(N__29683));
    InMux I__5113 (
            .O(N__29736),
            .I(N__29683));
    InMux I__5112 (
            .O(N__29735),
            .I(N__29683));
    InMux I__5111 (
            .O(N__29734),
            .I(N__29674));
    InMux I__5110 (
            .O(N__29733),
            .I(N__29674));
    InMux I__5109 (
            .O(N__29732),
            .I(N__29674));
    InMux I__5108 (
            .O(N__29731),
            .I(N__29674));
    Span4Mux_v I__5107 (
            .O(N__29728),
            .I(N__29667));
    LocalMux I__5106 (
            .O(N__29719),
            .I(N__29667));
    LocalMux I__5105 (
            .O(N__29710),
            .I(N__29667));
    InMux I__5104 (
            .O(N__29709),
            .I(N__29658));
    InMux I__5103 (
            .O(N__29708),
            .I(N__29658));
    InMux I__5102 (
            .O(N__29707),
            .I(N__29658));
    InMux I__5101 (
            .O(N__29706),
            .I(N__29658));
    LocalMux I__5100 (
            .O(N__29701),
            .I(N__29645));
    LocalMux I__5099 (
            .O(N__29692),
            .I(N__29645));
    LocalMux I__5098 (
            .O(N__29683),
            .I(N__29645));
    LocalMux I__5097 (
            .O(N__29674),
            .I(N__29645));
    Span4Mux_h I__5096 (
            .O(N__29667),
            .I(N__29645));
    LocalMux I__5095 (
            .O(N__29658),
            .I(N__29645));
    Span4Mux_v I__5094 (
            .O(N__29645),
            .I(N__29642));
    Odrv4 I__5093 (
            .O(N__29642),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    CascadeMux I__5092 (
            .O(N__29639),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    InMux I__5091 (
            .O(N__29636),
            .I(N__29633));
    LocalMux I__5090 (
            .O(N__29633),
            .I(N__29629));
    InMux I__5089 (
            .O(N__29632),
            .I(N__29626));
    Span4Mux_v I__5088 (
            .O(N__29629),
            .I(N__29623));
    LocalMux I__5087 (
            .O(N__29626),
            .I(N__29620));
    Sp12to4 I__5086 (
            .O(N__29623),
            .I(N__29617));
    Span4Mux_h I__5085 (
            .O(N__29620),
            .I(N__29614));
    Span12Mux_s11_h I__5084 (
            .O(N__29617),
            .I(N__29611));
    Odrv4 I__5083 (
            .O(N__29614),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv12 I__5082 (
            .O(N__29611),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__5081 (
            .O(N__29606),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__5080 (
            .O(N__29603),
            .I(bfn_11_14_0_));
    InMux I__5079 (
            .O(N__29600),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__5078 (
            .O(N__29597),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__5077 (
            .O(N__29594),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__5076 (
            .O(N__29591),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__5075 (
            .O(N__29588),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__5074 (
            .O(N__29585),
            .I(N__29581));
    InMux I__5073 (
            .O(N__29584),
            .I(N__29578));
    LocalMux I__5072 (
            .O(N__29581),
            .I(N__29572));
    LocalMux I__5071 (
            .O(N__29578),
            .I(N__29572));
    InMux I__5070 (
            .O(N__29577),
            .I(N__29567));
    Span4Mux_v I__5069 (
            .O(N__29572),
            .I(N__29564));
    InMux I__5068 (
            .O(N__29571),
            .I(N__29559));
    InMux I__5067 (
            .O(N__29570),
            .I(N__29559));
    LocalMux I__5066 (
            .O(N__29567),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__5065 (
            .O(N__29564),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__5064 (
            .O(N__29559),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__5063 (
            .O(N__29552),
            .I(N__29549));
    LocalMux I__5062 (
            .O(N__29549),
            .I(N__29545));
    InMux I__5061 (
            .O(N__29548),
            .I(N__29541));
    Span4Mux_v I__5060 (
            .O(N__29545),
            .I(N__29538));
    InMux I__5059 (
            .O(N__29544),
            .I(N__29535));
    LocalMux I__5058 (
            .O(N__29541),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__5057 (
            .O(N__29538),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    LocalMux I__5056 (
            .O(N__29535),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__5055 (
            .O(N__29528),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__5054 (
            .O(N__29525),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__5053 (
            .O(N__29522),
            .I(bfn_11_13_0_));
    InMux I__5052 (
            .O(N__29519),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__5051 (
            .O(N__29516),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__5050 (
            .O(N__29513),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__5049 (
            .O(N__29510),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__5048 (
            .O(N__29507),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__5047 (
            .O(N__29504),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__5046 (
            .O(N__29501),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__5045 (
            .O(N__29498),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__5044 (
            .O(N__29495),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__5043 (
            .O(N__29492),
            .I(bfn_11_12_0_));
    InMux I__5042 (
            .O(N__29489),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__5041 (
            .O(N__29486),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__5040 (
            .O(N__29483),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__5039 (
            .O(N__29480),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__5038 (
            .O(N__29477),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    CascadeMux I__5037 (
            .O(N__29474),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ));
    InMux I__5036 (
            .O(N__29471),
            .I(N__29465));
    InMux I__5035 (
            .O(N__29470),
            .I(N__29465));
    LocalMux I__5034 (
            .O(N__29465),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__5033 (
            .O(N__29462),
            .I(N__29459));
    LocalMux I__5032 (
            .O(N__29459),
            .I(N__29456));
    Span4Mux_v I__5031 (
            .O(N__29456),
            .I(N__29450));
    InMux I__5030 (
            .O(N__29455),
            .I(N__29443));
    InMux I__5029 (
            .O(N__29454),
            .I(N__29443));
    InMux I__5028 (
            .O(N__29453),
            .I(N__29443));
    Odrv4 I__5027 (
            .O(N__29450),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__5026 (
            .O(N__29443),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__5025 (
            .O(N__29438),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__5024 (
            .O(N__29435),
            .I(bfn_11_11_0_));
    InMux I__5023 (
            .O(N__29432),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__5022 (
            .O(N__29429),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__5021 (
            .O(N__29426),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__5020 (
            .O(N__29423),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__5019 (
            .O(N__29420),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__5018 (
            .O(N__29417),
            .I(N__29413));
    InMux I__5017 (
            .O(N__29416),
            .I(N__29409));
    LocalMux I__5016 (
            .O(N__29413),
            .I(N__29406));
    InMux I__5015 (
            .O(N__29412),
            .I(N__29403));
    LocalMux I__5014 (
            .O(N__29409),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    Odrv4 I__5013 (
            .O(N__29406),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__5012 (
            .O(N__29403),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__5011 (
            .O(N__29396),
            .I(N__29393));
    LocalMux I__5010 (
            .O(N__29393),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    CascadeMux I__5009 (
            .O(N__29390),
            .I(N__29387));
    InMux I__5008 (
            .O(N__29387),
            .I(N__29384));
    LocalMux I__5007 (
            .O(N__29384),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    InMux I__5006 (
            .O(N__29381),
            .I(N__29378));
    LocalMux I__5005 (
            .O(N__29378),
            .I(N__29375));
    Span4Mux_h I__5004 (
            .O(N__29375),
            .I(N__29371));
    InMux I__5003 (
            .O(N__29374),
            .I(N__29368));
    Odrv4 I__5002 (
            .O(N__29371),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    LocalMux I__5001 (
            .O(N__29368),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    CascadeMux I__5000 (
            .O(N__29363),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17_cascade_));
    CascadeMux I__4999 (
            .O(N__29360),
            .I(N__29357));
    InMux I__4998 (
            .O(N__29357),
            .I(N__29351));
    InMux I__4997 (
            .O(N__29356),
            .I(N__29351));
    LocalMux I__4996 (
            .O(N__29351),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__4995 (
            .O(N__29348),
            .I(N__29345));
    LocalMux I__4994 (
            .O(N__29345),
            .I(N__29341));
    InMux I__4993 (
            .O(N__29344),
            .I(N__29337));
    Span4Mux_h I__4992 (
            .O(N__29341),
            .I(N__29334));
    InMux I__4991 (
            .O(N__29340),
            .I(N__29331));
    LocalMux I__4990 (
            .O(N__29337),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    Odrv4 I__4989 (
            .O(N__29334),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    LocalMux I__4988 (
            .O(N__29331),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__4987 (
            .O(N__29324),
            .I(N__29318));
    InMux I__4986 (
            .O(N__29323),
            .I(N__29318));
    LocalMux I__4985 (
            .O(N__29318),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__4984 (
            .O(N__29315),
            .I(N__29311));
    InMux I__4983 (
            .O(N__29314),
            .I(N__29308));
    InMux I__4982 (
            .O(N__29311),
            .I(N__29304));
    LocalMux I__4981 (
            .O(N__29308),
            .I(N__29301));
    InMux I__4980 (
            .O(N__29307),
            .I(N__29298));
    LocalMux I__4979 (
            .O(N__29304),
            .I(N__29293));
    Span4Mux_h I__4978 (
            .O(N__29301),
            .I(N__29293));
    LocalMux I__4977 (
            .O(N__29298),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    Odrv4 I__4976 (
            .O(N__29293),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__4975 (
            .O(N__29288),
            .I(N__29285));
    LocalMux I__4974 (
            .O(N__29285),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__4973 (
            .O(N__29282),
            .I(N__29279));
    LocalMux I__4972 (
            .O(N__29279),
            .I(N__29276));
    Odrv12 I__4971 (
            .O(N__29276),
            .I(\phase_controller_inst1.N_49_0 ));
    InMux I__4970 (
            .O(N__29273),
            .I(N__29267));
    InMux I__4969 (
            .O(N__29272),
            .I(N__29264));
    InMux I__4968 (
            .O(N__29271),
            .I(N__29259));
    InMux I__4967 (
            .O(N__29270),
            .I(N__29259));
    LocalMux I__4966 (
            .O(N__29267),
            .I(N__29254));
    LocalMux I__4965 (
            .O(N__29264),
            .I(N__29254));
    LocalMux I__4964 (
            .O(N__29259),
            .I(N__29251));
    Span4Mux_v I__4963 (
            .O(N__29254),
            .I(N__29248));
    Span4Mux_h I__4962 (
            .O(N__29251),
            .I(N__29245));
    Odrv4 I__4961 (
            .O(N__29248),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv4 I__4960 (
            .O(N__29245),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__4959 (
            .O(N__29240),
            .I(N__29236));
    InMux I__4958 (
            .O(N__29239),
            .I(N__29233));
    LocalMux I__4957 (
            .O(N__29236),
            .I(N__29230));
    LocalMux I__4956 (
            .O(N__29233),
            .I(N__29225));
    Span4Mux_v I__4955 (
            .O(N__29230),
            .I(N__29222));
    InMux I__4954 (
            .O(N__29229),
            .I(N__29219));
    InMux I__4953 (
            .O(N__29228),
            .I(N__29216));
    Span4Mux_h I__4952 (
            .O(N__29225),
            .I(N__29213));
    Odrv4 I__4951 (
            .O(N__29222),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__4950 (
            .O(N__29219),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__4949 (
            .O(N__29216),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv4 I__4948 (
            .O(N__29213),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__4947 (
            .O(N__29204),
            .I(N__29201));
    LocalMux I__4946 (
            .O(N__29201),
            .I(N__29197));
    InMux I__4945 (
            .O(N__29200),
            .I(N__29193));
    Span4Mux_h I__4944 (
            .O(N__29197),
            .I(N__29190));
    InMux I__4943 (
            .O(N__29196),
            .I(N__29187));
    LocalMux I__4942 (
            .O(N__29193),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv4 I__4941 (
            .O(N__29190),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    LocalMux I__4940 (
            .O(N__29187),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__4939 (
            .O(N__29180),
            .I(N__29176));
    InMux I__4938 (
            .O(N__29179),
            .I(N__29172));
    LocalMux I__4937 (
            .O(N__29176),
            .I(N__29169));
    InMux I__4936 (
            .O(N__29175),
            .I(N__29166));
    LocalMux I__4935 (
            .O(N__29172),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv4 I__4934 (
            .O(N__29169),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    LocalMux I__4933 (
            .O(N__29166),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    CascadeMux I__4932 (
            .O(N__29159),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ));
    InMux I__4931 (
            .O(N__29156),
            .I(N__29153));
    LocalMux I__4930 (
            .O(N__29153),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ));
    InMux I__4929 (
            .O(N__29150),
            .I(N__29147));
    LocalMux I__4928 (
            .O(N__29147),
            .I(N__29144));
    Odrv12 I__4927 (
            .O(N__29144),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ));
    InMux I__4926 (
            .O(N__29141),
            .I(N__29138));
    LocalMux I__4925 (
            .O(N__29138),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ));
    CascadeMux I__4924 (
            .O(N__29135),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ));
    InMux I__4923 (
            .O(N__29132),
            .I(N__29129));
    LocalMux I__4922 (
            .O(N__29129),
            .I(\phase_controller_inst2.N_51_0 ));
    InMux I__4921 (
            .O(N__29126),
            .I(N__29123));
    LocalMux I__4920 (
            .O(N__29123),
            .I(N__29120));
    Span4Mux_h I__4919 (
            .O(N__29120),
            .I(N__29114));
    InMux I__4918 (
            .O(N__29119),
            .I(N__29111));
    InMux I__4917 (
            .O(N__29118),
            .I(N__29108));
    CascadeMux I__4916 (
            .O(N__29117),
            .I(N__29105));
    Sp12to4 I__4915 (
            .O(N__29114),
            .I(N__29098));
    LocalMux I__4914 (
            .O(N__29111),
            .I(N__29098));
    LocalMux I__4913 (
            .O(N__29108),
            .I(N__29098));
    InMux I__4912 (
            .O(N__29105),
            .I(N__29095));
    Span12Mux_v I__4911 (
            .O(N__29098),
            .I(N__29092));
    LocalMux I__4910 (
            .O(N__29095),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv12 I__4909 (
            .O(N__29092),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__4908 (
            .O(N__29087),
            .I(N__29080));
    InMux I__4907 (
            .O(N__29086),
            .I(N__29080));
    InMux I__4906 (
            .O(N__29085),
            .I(N__29077));
    LocalMux I__4905 (
            .O(N__29080),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__4904 (
            .O(N__29077),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__4903 (
            .O(N__29072),
            .I(N__29069));
    InMux I__4902 (
            .O(N__29069),
            .I(N__29065));
    InMux I__4901 (
            .O(N__29068),
            .I(N__29062));
    LocalMux I__4900 (
            .O(N__29065),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__4899 (
            .O(N__29062),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__4898 (
            .O(N__29057),
            .I(N__29054));
    LocalMux I__4897 (
            .O(N__29054),
            .I(N__29051));
    Odrv12 I__4896 (
            .O(N__29051),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    InMux I__4895 (
            .O(N__29048),
            .I(N__29045));
    LocalMux I__4894 (
            .O(N__29045),
            .I(N__29042));
    Odrv12 I__4893 (
            .O(N__29042),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ));
    InMux I__4892 (
            .O(N__29039),
            .I(N__29036));
    LocalMux I__4891 (
            .O(N__29036),
            .I(N__29033));
    Odrv12 I__4890 (
            .O(N__29033),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ));
    InMux I__4889 (
            .O(N__29030),
            .I(N__29027));
    LocalMux I__4888 (
            .O(N__29027),
            .I(N__29024));
    Odrv12 I__4887 (
            .O(N__29024),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ));
    InMux I__4886 (
            .O(N__29021),
            .I(N__29016));
    InMux I__4885 (
            .O(N__29020),
            .I(N__29012));
    InMux I__4884 (
            .O(N__29019),
            .I(N__29009));
    LocalMux I__4883 (
            .O(N__29016),
            .I(N__29006));
    InMux I__4882 (
            .O(N__29015),
            .I(N__29003));
    LocalMux I__4881 (
            .O(N__29012),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__4880 (
            .O(N__29009),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv12 I__4879 (
            .O(N__29006),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__4878 (
            .O(N__29003),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    IoInMux I__4877 (
            .O(N__28994),
            .I(N__28991));
    LocalMux I__4876 (
            .O(N__28991),
            .I(N__28988));
    IoSpan4Mux I__4875 (
            .O(N__28988),
            .I(N__28985));
    Span4Mux_s3_v I__4874 (
            .O(N__28985),
            .I(N__28982));
    Span4Mux_v I__4873 (
            .O(N__28982),
            .I(N__28979));
    Odrv4 I__4872 (
            .O(N__28979),
            .I(s4_phy_c));
    InMux I__4871 (
            .O(N__28976),
            .I(N__28971));
    InMux I__4870 (
            .O(N__28975),
            .I(N__28968));
    InMux I__4869 (
            .O(N__28974),
            .I(N__28965));
    LocalMux I__4868 (
            .O(N__28971),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__4867 (
            .O(N__28968),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__4866 (
            .O(N__28965),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__4865 (
            .O(N__28958),
            .I(N__28954));
    InMux I__4864 (
            .O(N__28957),
            .I(N__28950));
    LocalMux I__4863 (
            .O(N__28954),
            .I(N__28947));
    InMux I__4862 (
            .O(N__28953),
            .I(N__28944));
    LocalMux I__4861 (
            .O(N__28950),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv4 I__4860 (
            .O(N__28947),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    LocalMux I__4859 (
            .O(N__28944),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    InMux I__4858 (
            .O(N__28937),
            .I(N__28933));
    InMux I__4857 (
            .O(N__28936),
            .I(N__28930));
    LocalMux I__4856 (
            .O(N__28933),
            .I(N__28927));
    LocalMux I__4855 (
            .O(N__28930),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    Odrv4 I__4854 (
            .O(N__28927),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    CEMux I__4853 (
            .O(N__28922),
            .I(N__28889));
    CEMux I__4852 (
            .O(N__28921),
            .I(N__28889));
    CEMux I__4851 (
            .O(N__28920),
            .I(N__28889));
    CEMux I__4850 (
            .O(N__28919),
            .I(N__28889));
    CEMux I__4849 (
            .O(N__28918),
            .I(N__28889));
    CEMux I__4848 (
            .O(N__28917),
            .I(N__28889));
    CEMux I__4847 (
            .O(N__28916),
            .I(N__28889));
    CEMux I__4846 (
            .O(N__28915),
            .I(N__28889));
    CEMux I__4845 (
            .O(N__28914),
            .I(N__28889));
    CEMux I__4844 (
            .O(N__28913),
            .I(N__28889));
    CEMux I__4843 (
            .O(N__28912),
            .I(N__28889));
    GlobalMux I__4842 (
            .O(N__28889),
            .I(N__28886));
    gio2CtrlBuf I__4841 (
            .O(N__28886),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    InMux I__4840 (
            .O(N__28883),
            .I(N__28878));
    InMux I__4839 (
            .O(N__28882),
            .I(N__28873));
    InMux I__4838 (
            .O(N__28881),
            .I(N__28873));
    LocalMux I__4837 (
            .O(N__28878),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__4836 (
            .O(N__28873),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    CascadeMux I__4835 (
            .O(N__28868),
            .I(N__28863));
    InMux I__4834 (
            .O(N__28867),
            .I(N__28857));
    InMux I__4833 (
            .O(N__28866),
            .I(N__28857));
    InMux I__4832 (
            .O(N__28863),
            .I(N__28852));
    InMux I__4831 (
            .O(N__28862),
            .I(N__28852));
    LocalMux I__4830 (
            .O(N__28857),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__4829 (
            .O(N__28852),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__4828 (
            .O(N__28847),
            .I(N__28844));
    LocalMux I__4827 (
            .O(N__28844),
            .I(\phase_controller_inst2.test_0_sqmuxa ));
    InMux I__4826 (
            .O(N__28841),
            .I(N__28838));
    LocalMux I__4825 (
            .O(N__28838),
            .I(N__28835));
    Span4Mux_v I__4824 (
            .O(N__28835),
            .I(N__28831));
    InMux I__4823 (
            .O(N__28834),
            .I(N__28828));
    Span4Mux_h I__4822 (
            .O(N__28831),
            .I(N__28825));
    LocalMux I__4821 (
            .O(N__28828),
            .I(N__28822));
    Span4Mux_v I__4820 (
            .O(N__28825),
            .I(N__28816));
    Span4Mux_v I__4819 (
            .O(N__28822),
            .I(N__28813));
    InMux I__4818 (
            .O(N__28821),
            .I(N__28808));
    InMux I__4817 (
            .O(N__28820),
            .I(N__28808));
    InMux I__4816 (
            .O(N__28819),
            .I(N__28805));
    Span4Mux_v I__4815 (
            .O(N__28816),
            .I(N__28802));
    Span4Mux_v I__4814 (
            .O(N__28813),
            .I(N__28795));
    LocalMux I__4813 (
            .O(N__28808),
            .I(N__28795));
    LocalMux I__4812 (
            .O(N__28805),
            .I(N__28795));
    Odrv4 I__4811 (
            .O(N__28802),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__4810 (
            .O(N__28795),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    CascadeMux I__4809 (
            .O(N__28790),
            .I(N__28787));
    InMux I__4808 (
            .O(N__28787),
            .I(N__28784));
    LocalMux I__4807 (
            .O(N__28784),
            .I(N__28780));
    InMux I__4806 (
            .O(N__28783),
            .I(N__28777));
    Span4Mux_v I__4805 (
            .O(N__28780),
            .I(N__28774));
    LocalMux I__4804 (
            .O(N__28777),
            .I(N__28771));
    Span4Mux_h I__4803 (
            .O(N__28774),
            .I(N__28768));
    Span12Mux_s11_v I__4802 (
            .O(N__28771),
            .I(N__28763));
    Span4Mux_v I__4801 (
            .O(N__28768),
            .I(N__28760));
    InMux I__4800 (
            .O(N__28767),
            .I(N__28755));
    InMux I__4799 (
            .O(N__28766),
            .I(N__28755));
    Odrv12 I__4798 (
            .O(N__28763),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__4797 (
            .O(N__28760),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__4796 (
            .O(N__28755),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__4795 (
            .O(N__28748),
            .I(N__28744));
    InMux I__4794 (
            .O(N__28747),
            .I(N__28740));
    LocalMux I__4793 (
            .O(N__28744),
            .I(N__28737));
    InMux I__4792 (
            .O(N__28743),
            .I(N__28734));
    LocalMux I__4791 (
            .O(N__28740),
            .I(N__28731));
    Span4Mux_h I__4790 (
            .O(N__28737),
            .I(N__28728));
    LocalMux I__4789 (
            .O(N__28734),
            .I(N__28725));
    Span4Mux_v I__4788 (
            .O(N__28731),
            .I(N__28720));
    Span4Mux_v I__4787 (
            .O(N__28728),
            .I(N__28720));
    Span4Mux_h I__4786 (
            .O(N__28725),
            .I(N__28717));
    Odrv4 I__4785 (
            .O(N__28720),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__4784 (
            .O(N__28717),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__4783 (
            .O(N__28712),
            .I(N__28706));
    InMux I__4782 (
            .O(N__28711),
            .I(N__28706));
    LocalMux I__4781 (
            .O(N__28706),
            .I(N__28703));
    Span4Mux_v I__4780 (
            .O(N__28703),
            .I(N__28699));
    InMux I__4779 (
            .O(N__28702),
            .I(N__28696));
    Span4Mux_h I__4778 (
            .O(N__28699),
            .I(N__28693));
    LocalMux I__4777 (
            .O(N__28696),
            .I(N__28690));
    Sp12to4 I__4776 (
            .O(N__28693),
            .I(N__28685));
    Span12Mux_h I__4775 (
            .O(N__28690),
            .I(N__28685));
    Span12Mux_v I__4774 (
            .O(N__28685),
            .I(N__28682));
    Odrv12 I__4773 (
            .O(N__28682),
            .I(il_min_comp2_c));
    InMux I__4772 (
            .O(N__28679),
            .I(N__28675));
    InMux I__4771 (
            .O(N__28678),
            .I(N__28672));
    LocalMux I__4770 (
            .O(N__28675),
            .I(\phase_controller_inst2.N_58 ));
    LocalMux I__4769 (
            .O(N__28672),
            .I(\phase_controller_inst2.N_58 ));
    InMux I__4768 (
            .O(N__28667),
            .I(N__28663));
    InMux I__4767 (
            .O(N__28666),
            .I(N__28660));
    LocalMux I__4766 (
            .O(N__28663),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    LocalMux I__4765 (
            .O(N__28660),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    InMux I__4764 (
            .O(N__28655),
            .I(N__28651));
    InMux I__4763 (
            .O(N__28654),
            .I(N__28648));
    LocalMux I__4762 (
            .O(N__28651),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    LocalMux I__4761 (
            .O(N__28648),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    InMux I__4760 (
            .O(N__28643),
            .I(N__28640));
    LocalMux I__4759 (
            .O(N__28640),
            .I(N__28635));
    InMux I__4758 (
            .O(N__28639),
            .I(N__28632));
    InMux I__4757 (
            .O(N__28638),
            .I(N__28629));
    Span4Mux_h I__4756 (
            .O(N__28635),
            .I(N__28626));
    LocalMux I__4755 (
            .O(N__28632),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    LocalMux I__4754 (
            .O(N__28629),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    Odrv4 I__4753 (
            .O(N__28626),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    CascadeMux I__4752 (
            .O(N__28619),
            .I(N__28616));
    InMux I__4751 (
            .O(N__28616),
            .I(N__28613));
    LocalMux I__4750 (
            .O(N__28613),
            .I(N__28610));
    Odrv12 I__4749 (
            .O(N__28610),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__4748 (
            .O(N__28607),
            .I(N__28604));
    LocalMux I__4747 (
            .O(N__28604),
            .I(N__28601));
    Odrv12 I__4746 (
            .O(N__28601),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__4745 (
            .O(N__28598),
            .I(N__28595));
    LocalMux I__4744 (
            .O(N__28595),
            .I(N__28592));
    Odrv12 I__4743 (
            .O(N__28592),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__4742 (
            .O(N__28589),
            .I(N__28586));
    LocalMux I__4741 (
            .O(N__28586),
            .I(N__28583));
    Span4Mux_h I__4740 (
            .O(N__28583),
            .I(N__28579));
    InMux I__4739 (
            .O(N__28582),
            .I(N__28575));
    Sp12to4 I__4738 (
            .O(N__28579),
            .I(N__28572));
    InMux I__4737 (
            .O(N__28578),
            .I(N__28569));
    LocalMux I__4736 (
            .O(N__28575),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv12 I__4735 (
            .O(N__28572),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    LocalMux I__4734 (
            .O(N__28569),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__4733 (
            .O(N__28562),
            .I(N__28557));
    InMux I__4732 (
            .O(N__28561),
            .I(N__28554));
    InMux I__4731 (
            .O(N__28560),
            .I(N__28551));
    LocalMux I__4730 (
            .O(N__28557),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    LocalMux I__4729 (
            .O(N__28554),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    LocalMux I__4728 (
            .O(N__28551),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    InMux I__4727 (
            .O(N__28544),
            .I(N__28538));
    InMux I__4726 (
            .O(N__28543),
            .I(N__28538));
    LocalMux I__4725 (
            .O(N__28538),
            .I(N__28535));
    Span4Mux_v I__4724 (
            .O(N__28535),
            .I(N__28532));
    Odrv4 I__4723 (
            .O(N__28532),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    InMux I__4722 (
            .O(N__28529),
            .I(N__28523));
    InMux I__4721 (
            .O(N__28528),
            .I(N__28523));
    LocalMux I__4720 (
            .O(N__28523),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    CascadeMux I__4719 (
            .O(N__28520),
            .I(N__28517));
    InMux I__4718 (
            .O(N__28517),
            .I(N__28514));
    LocalMux I__4717 (
            .O(N__28514),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    InMux I__4716 (
            .O(N__28511),
            .I(N__28508));
    LocalMux I__4715 (
            .O(N__28508),
            .I(N__28503));
    InMux I__4714 (
            .O(N__28507),
            .I(N__28500));
    InMux I__4713 (
            .O(N__28506),
            .I(N__28497));
    Span4Mux_v I__4712 (
            .O(N__28503),
            .I(N__28494));
    LocalMux I__4711 (
            .O(N__28500),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    LocalMux I__4710 (
            .O(N__28497),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv4 I__4709 (
            .O(N__28494),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__4708 (
            .O(N__28487),
            .I(N__28484));
    LocalMux I__4707 (
            .O(N__28484),
            .I(N__28481));
    Odrv12 I__4706 (
            .O(N__28481),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__4705 (
            .O(N__28478),
            .I(N__28475));
    LocalMux I__4704 (
            .O(N__28475),
            .I(N__28472));
    Span4Mux_h I__4703 (
            .O(N__28472),
            .I(N__28468));
    InMux I__4702 (
            .O(N__28471),
            .I(N__28465));
    Odrv4 I__4701 (
            .O(N__28468),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    LocalMux I__4700 (
            .O(N__28465),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__4699 (
            .O(N__28460),
            .I(N__28457));
    LocalMux I__4698 (
            .O(N__28457),
            .I(N__28454));
    Span4Mux_v I__4697 (
            .O(N__28454),
            .I(N__28451));
    Odrv4 I__4696 (
            .O(N__28451),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__4695 (
            .O(N__28448),
            .I(N__28445));
    InMux I__4694 (
            .O(N__28445),
            .I(N__28442));
    LocalMux I__4693 (
            .O(N__28442),
            .I(N__28439));
    Odrv4 I__4692 (
            .O(N__28439),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    InMux I__4691 (
            .O(N__28436),
            .I(N__28433));
    LocalMux I__4690 (
            .O(N__28433),
            .I(N__28430));
    Odrv4 I__4689 (
            .O(N__28430),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    InMux I__4688 (
            .O(N__28427),
            .I(N__28424));
    LocalMux I__4687 (
            .O(N__28424),
            .I(N__28421));
    Span4Mux_h I__4686 (
            .O(N__28421),
            .I(N__28417));
    InMux I__4685 (
            .O(N__28420),
            .I(N__28414));
    Odrv4 I__4684 (
            .O(N__28417),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    LocalMux I__4683 (
            .O(N__28414),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    CascadeMux I__4682 (
            .O(N__28409),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29_cascade_));
    CascadeMux I__4681 (
            .O(N__28406),
            .I(N__28403));
    InMux I__4680 (
            .O(N__28403),
            .I(N__28397));
    InMux I__4679 (
            .O(N__28402),
            .I(N__28397));
    LocalMux I__4678 (
            .O(N__28397),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    InMux I__4677 (
            .O(N__28394),
            .I(N__28389));
    InMux I__4676 (
            .O(N__28393),
            .I(N__28386));
    InMux I__4675 (
            .O(N__28392),
            .I(N__28383));
    LocalMux I__4674 (
            .O(N__28389),
            .I(N__28380));
    LocalMux I__4673 (
            .O(N__28386),
            .I(N__28377));
    LocalMux I__4672 (
            .O(N__28383),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv12 I__4671 (
            .O(N__28380),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv4 I__4670 (
            .O(N__28377),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__4669 (
            .O(N__28370),
            .I(N__28364));
    InMux I__4668 (
            .O(N__28369),
            .I(N__28364));
    LocalMux I__4667 (
            .O(N__28364),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    InMux I__4666 (
            .O(N__28361),
            .I(N__28358));
    LocalMux I__4665 (
            .O(N__28358),
            .I(N__28355));
    Odrv4 I__4664 (
            .O(N__28355),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    InMux I__4663 (
            .O(N__28352),
            .I(N__28349));
    LocalMux I__4662 (
            .O(N__28349),
            .I(N__28346));
    Odrv12 I__4661 (
            .O(N__28346),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    CascadeMux I__4660 (
            .O(N__28343),
            .I(N__28340));
    InMux I__4659 (
            .O(N__28340),
            .I(N__28337));
    LocalMux I__4658 (
            .O(N__28337),
            .I(N__28334));
    Span4Mux_v I__4657 (
            .O(N__28334),
            .I(N__28331));
    Odrv4 I__4656 (
            .O(N__28331),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    InMux I__4655 (
            .O(N__28328),
            .I(N__28325));
    LocalMux I__4654 (
            .O(N__28325),
            .I(N__28322));
    Odrv4 I__4653 (
            .O(N__28322),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    CascadeMux I__4652 (
            .O(N__28319),
            .I(N__28316));
    InMux I__4651 (
            .O(N__28316),
            .I(N__28313));
    LocalMux I__4650 (
            .O(N__28313),
            .I(N__28310));
    Odrv4 I__4649 (
            .O(N__28310),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    CascadeMux I__4648 (
            .O(N__28307),
            .I(N__28304));
    InMux I__4647 (
            .O(N__28304),
            .I(N__28301));
    LocalMux I__4646 (
            .O(N__28301),
            .I(N__28298));
    Span4Mux_h I__4645 (
            .O(N__28298),
            .I(N__28295));
    Odrv4 I__4644 (
            .O(N__28295),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ));
    InMux I__4643 (
            .O(N__28292),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    InMux I__4642 (
            .O(N__28289),
            .I(N__28286));
    LocalMux I__4641 (
            .O(N__28286),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    CascadeMux I__4640 (
            .O(N__28283),
            .I(N__28280));
    InMux I__4639 (
            .O(N__28280),
            .I(N__28277));
    LocalMux I__4638 (
            .O(N__28277),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__4637 (
            .O(N__28274),
            .I(N__28271));
    LocalMux I__4636 (
            .O(N__28271),
            .I(N__28268));
    Span4Mux_h I__4635 (
            .O(N__28268),
            .I(N__28265));
    Odrv4 I__4634 (
            .O(N__28265),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__4633 (
            .O(N__28262),
            .I(N__28259));
    InMux I__4632 (
            .O(N__28259),
            .I(N__28256));
    LocalMux I__4631 (
            .O(N__28256),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__4630 (
            .O(N__28253),
            .I(N__28250));
    LocalMux I__4629 (
            .O(N__28250),
            .I(N__28247));
    Span4Mux_h I__4628 (
            .O(N__28247),
            .I(N__28244));
    Odrv4 I__4627 (
            .O(N__28244),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__4626 (
            .O(N__28241),
            .I(N__28238));
    InMux I__4625 (
            .O(N__28238),
            .I(N__28235));
    LocalMux I__4624 (
            .O(N__28235),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__4623 (
            .O(N__28232),
            .I(N__28229));
    InMux I__4622 (
            .O(N__28229),
            .I(N__28226));
    LocalMux I__4621 (
            .O(N__28226),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__4620 (
            .O(N__28223),
            .I(N__28220));
    InMux I__4619 (
            .O(N__28220),
            .I(N__28217));
    LocalMux I__4618 (
            .O(N__28217),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__4617 (
            .O(N__28214),
            .I(N__28211));
    InMux I__4616 (
            .O(N__28211),
            .I(N__28208));
    LocalMux I__4615 (
            .O(N__28208),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__4614 (
            .O(N__28205),
            .I(N__28202));
    LocalMux I__4613 (
            .O(N__28202),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__4612 (
            .O(N__28199),
            .I(N__28196));
    LocalMux I__4611 (
            .O(N__28196),
            .I(N__28193));
    Odrv12 I__4610 (
            .O(N__28193),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    CascadeMux I__4609 (
            .O(N__28190),
            .I(N__28187));
    InMux I__4608 (
            .O(N__28187),
            .I(N__28184));
    LocalMux I__4607 (
            .O(N__28184),
            .I(N__28181));
    Odrv12 I__4606 (
            .O(N__28181),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__4605 (
            .O(N__28178),
            .I(N__28175));
    LocalMux I__4604 (
            .O(N__28175),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    CascadeMux I__4603 (
            .O(N__28172),
            .I(N__28169));
    InMux I__4602 (
            .O(N__28169),
            .I(N__28166));
    LocalMux I__4601 (
            .O(N__28166),
            .I(N__28163));
    Odrv4 I__4600 (
            .O(N__28163),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    InMux I__4599 (
            .O(N__28160),
            .I(N__28157));
    LocalMux I__4598 (
            .O(N__28157),
            .I(N__28154));
    Odrv4 I__4597 (
            .O(N__28154),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__4596 (
            .O(N__28151),
            .I(N__28148));
    InMux I__4595 (
            .O(N__28148),
            .I(N__28145));
    LocalMux I__4594 (
            .O(N__28145),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__4593 (
            .O(N__28142),
            .I(N__28139));
    LocalMux I__4592 (
            .O(N__28139),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__4591 (
            .O(N__28136),
            .I(N__28133));
    InMux I__4590 (
            .O(N__28133),
            .I(N__28130));
    LocalMux I__4589 (
            .O(N__28130),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__4588 (
            .O(N__28127),
            .I(N__28124));
    LocalMux I__4587 (
            .O(N__28124),
            .I(N__28121));
    Odrv4 I__4586 (
            .O(N__28121),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__4585 (
            .O(N__28118),
            .I(N__28115));
    InMux I__4584 (
            .O(N__28115),
            .I(N__28112));
    LocalMux I__4583 (
            .O(N__28112),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__4582 (
            .O(N__28109),
            .I(N__28106));
    InMux I__4581 (
            .O(N__28106),
            .I(N__28103));
    LocalMux I__4580 (
            .O(N__28103),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__4579 (
            .O(N__28100),
            .I(N__28097));
    LocalMux I__4578 (
            .O(N__28097),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__4577 (
            .O(N__28094),
            .I(N__28091));
    InMux I__4576 (
            .O(N__28091),
            .I(N__28088));
    LocalMux I__4575 (
            .O(N__28088),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__4574 (
            .O(N__28085),
            .I(N__28082));
    InMux I__4573 (
            .O(N__28082),
            .I(N__28079));
    LocalMux I__4572 (
            .O(N__28079),
            .I(N__28076));
    Odrv4 I__4571 (
            .O(N__28076),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__4570 (
            .O(N__28073),
            .I(N__28070));
    LocalMux I__4569 (
            .O(N__28070),
            .I(N__28067));
    Odrv4 I__4568 (
            .O(N__28067),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__4567 (
            .O(N__28064),
            .I(N__28061));
    InMux I__4566 (
            .O(N__28061),
            .I(N__28058));
    LocalMux I__4565 (
            .O(N__28058),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__4564 (
            .O(N__28055),
            .I(N__28052));
    LocalMux I__4563 (
            .O(N__28052),
            .I(N__28049));
    Odrv4 I__4562 (
            .O(N__28049),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    InMux I__4561 (
            .O(N__28046),
            .I(N__28041));
    InMux I__4560 (
            .O(N__28045),
            .I(N__28038));
    InMux I__4559 (
            .O(N__28044),
            .I(N__28035));
    LocalMux I__4558 (
            .O(N__28041),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__4557 (
            .O(N__28038),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__4556 (
            .O(N__28035),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    InMux I__4555 (
            .O(N__28028),
            .I(N__28023));
    InMux I__4554 (
            .O(N__28027),
            .I(N__28020));
    InMux I__4553 (
            .O(N__28026),
            .I(N__28017));
    LocalMux I__4552 (
            .O(N__28023),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__4551 (
            .O(N__28020),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__4550 (
            .O(N__28017),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    InMux I__4549 (
            .O(N__28010),
            .I(N__28004));
    InMux I__4548 (
            .O(N__28009),
            .I(N__28004));
    LocalMux I__4547 (
            .O(N__28004),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    InMux I__4546 (
            .O(N__28001),
            .I(N__27997));
    InMux I__4545 (
            .O(N__28000),
            .I(N__27994));
    LocalMux I__4544 (
            .O(N__27997),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    LocalMux I__4543 (
            .O(N__27994),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    InMux I__4542 (
            .O(N__27989),
            .I(N__27984));
    InMux I__4541 (
            .O(N__27988),
            .I(N__27981));
    InMux I__4540 (
            .O(N__27987),
            .I(N__27978));
    LocalMux I__4539 (
            .O(N__27984),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    LocalMux I__4538 (
            .O(N__27981),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    LocalMux I__4537 (
            .O(N__27978),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    CascadeMux I__4536 (
            .O(N__27971),
            .I(N__27968));
    InMux I__4535 (
            .O(N__27968),
            .I(N__27965));
    LocalMux I__4534 (
            .O(N__27965),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__4533 (
            .O(N__27962),
            .I(N__27959));
    LocalMux I__4532 (
            .O(N__27959),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__4531 (
            .O(N__27956),
            .I(N__27953));
    LocalMux I__4530 (
            .O(N__27953),
            .I(N__27950));
    Odrv12 I__4529 (
            .O(N__27950),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ));
    InMux I__4528 (
            .O(N__27947),
            .I(N__27944));
    LocalMux I__4527 (
            .O(N__27944),
            .I(N__27941));
    Odrv12 I__4526 (
            .O(N__27941),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    IoInMux I__4525 (
            .O(N__27938),
            .I(N__27935));
    LocalMux I__4524 (
            .O(N__27935),
            .I(N__27932));
    Odrv12 I__4523 (
            .O(N__27932),
            .I(s3_phy_c));
    InMux I__4522 (
            .O(N__27929),
            .I(N__27926));
    LocalMux I__4521 (
            .O(N__27926),
            .I(N__27923));
    Glb2LocalMux I__4520 (
            .O(N__27923),
            .I(N__27920));
    GlobalMux I__4519 (
            .O(N__27920),
            .I(clk_12mhz));
    IoInMux I__4518 (
            .O(N__27917),
            .I(N__27914));
    LocalMux I__4517 (
            .O(N__27914),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__4516 (
            .O(N__27911),
            .I(N__27905));
    InMux I__4515 (
            .O(N__27910),
            .I(N__27905));
    LocalMux I__4514 (
            .O(N__27905),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__4513 (
            .O(N__27902),
            .I(N__27898));
    InMux I__4512 (
            .O(N__27901),
            .I(N__27893));
    InMux I__4511 (
            .O(N__27898),
            .I(N__27893));
    LocalMux I__4510 (
            .O(N__27893),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__4509 (
            .O(N__27890),
            .I(N__27886));
    InMux I__4508 (
            .O(N__27889),
            .I(N__27883));
    InMux I__4507 (
            .O(N__27886),
            .I(N__27879));
    LocalMux I__4506 (
            .O(N__27883),
            .I(N__27876));
    InMux I__4505 (
            .O(N__27882),
            .I(N__27873));
    LocalMux I__4504 (
            .O(N__27879),
            .I(N__27870));
    Span4Mux_h I__4503 (
            .O(N__27876),
            .I(N__27867));
    LocalMux I__4502 (
            .O(N__27873),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    Odrv12 I__4501 (
            .O(N__27870),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    Odrv4 I__4500 (
            .O(N__27867),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    InMux I__4499 (
            .O(N__27860),
            .I(N__27855));
    InMux I__4498 (
            .O(N__27859),
            .I(N__27852));
    InMux I__4497 (
            .O(N__27858),
            .I(N__27849));
    LocalMux I__4496 (
            .O(N__27855),
            .I(N__27844));
    LocalMux I__4495 (
            .O(N__27852),
            .I(N__27844));
    LocalMux I__4494 (
            .O(N__27849),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    Odrv4 I__4493 (
            .O(N__27844),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    CascadeMux I__4492 (
            .O(N__27839),
            .I(N__27836));
    InMux I__4491 (
            .O(N__27836),
            .I(N__27833));
    LocalMux I__4490 (
            .O(N__27833),
            .I(N__27830));
    Odrv12 I__4489 (
            .O(N__27830),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__4488 (
            .O(N__27827),
            .I(N__27824));
    LocalMux I__4487 (
            .O(N__27824),
            .I(N__27821));
    Odrv12 I__4486 (
            .O(N__27821),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    InMux I__4485 (
            .O(N__27818),
            .I(N__27815));
    LocalMux I__4484 (
            .O(N__27815),
            .I(N__27812));
    Odrv12 I__4483 (
            .O(N__27812),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    CascadeMux I__4482 (
            .O(N__27809),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_));
    CascadeMux I__4481 (
            .O(N__27806),
            .I(N__27803));
    InMux I__4480 (
            .O(N__27803),
            .I(N__27797));
    InMux I__4479 (
            .O(N__27802),
            .I(N__27797));
    LocalMux I__4478 (
            .O(N__27797),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    InMux I__4477 (
            .O(N__27794),
            .I(N__27788));
    InMux I__4476 (
            .O(N__27793),
            .I(N__27788));
    LocalMux I__4475 (
            .O(N__27788),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    InMux I__4474 (
            .O(N__27785),
            .I(N__27781));
    InMux I__4473 (
            .O(N__27784),
            .I(N__27778));
    LocalMux I__4472 (
            .O(N__27781),
            .I(N__27774));
    LocalMux I__4471 (
            .O(N__27778),
            .I(N__27771));
    InMux I__4470 (
            .O(N__27777),
            .I(N__27768));
    Span4Mux_h I__4469 (
            .O(N__27774),
            .I(N__27763));
    Span4Mux_v I__4468 (
            .O(N__27771),
            .I(N__27763));
    LocalMux I__4467 (
            .O(N__27768),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__4466 (
            .O(N__27763),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    CascadeMux I__4465 (
            .O(N__27758),
            .I(N__27754));
    CascadeMux I__4464 (
            .O(N__27757),
            .I(N__27751));
    InMux I__4463 (
            .O(N__27754),
            .I(N__27748));
    InMux I__4462 (
            .O(N__27751),
            .I(N__27745));
    LocalMux I__4461 (
            .O(N__27748),
            .I(N__27741));
    LocalMux I__4460 (
            .O(N__27745),
            .I(N__27738));
    InMux I__4459 (
            .O(N__27744),
            .I(N__27735));
    Span4Mux_h I__4458 (
            .O(N__27741),
            .I(N__27732));
    Span4Mux_v I__4457 (
            .O(N__27738),
            .I(N__27729));
    LocalMux I__4456 (
            .O(N__27735),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__4455 (
            .O(N__27732),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__4454 (
            .O(N__27729),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    CascadeMux I__4453 (
            .O(N__27722),
            .I(N__27719));
    InMux I__4452 (
            .O(N__27719),
            .I(N__27716));
    LocalMux I__4451 (
            .O(N__27716),
            .I(N__27713));
    Odrv4 I__4450 (
            .O(N__27713),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    InMux I__4449 (
            .O(N__27710),
            .I(N__27706));
    InMux I__4448 (
            .O(N__27709),
            .I(N__27703));
    LocalMux I__4447 (
            .O(N__27706),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    LocalMux I__4446 (
            .O(N__27703),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    InMux I__4445 (
            .O(N__27698),
            .I(N__27695));
    LocalMux I__4444 (
            .O(N__27695),
            .I(N__27691));
    InMux I__4443 (
            .O(N__27694),
            .I(N__27688));
    Odrv4 I__4442 (
            .O(N__27691),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    LocalMux I__4441 (
            .O(N__27688),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    InMux I__4440 (
            .O(N__27683),
            .I(N__27680));
    LocalMux I__4439 (
            .O(N__27680),
            .I(N__27676));
    InMux I__4438 (
            .O(N__27679),
            .I(N__27673));
    Odrv12 I__4437 (
            .O(N__27676),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    LocalMux I__4436 (
            .O(N__27673),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    InMux I__4435 (
            .O(N__27668),
            .I(N__27665));
    LocalMux I__4434 (
            .O(N__27665),
            .I(N__27661));
    InMux I__4433 (
            .O(N__27664),
            .I(N__27657));
    Span4Mux_v I__4432 (
            .O(N__27661),
            .I(N__27654));
    InMux I__4431 (
            .O(N__27660),
            .I(N__27651));
    LocalMux I__4430 (
            .O(N__27657),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    Odrv4 I__4429 (
            .O(N__27654),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__4428 (
            .O(N__27651),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    InMux I__4427 (
            .O(N__27644),
            .I(N__27641));
    LocalMux I__4426 (
            .O(N__27641),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    InMux I__4425 (
            .O(N__27638),
            .I(N__27635));
    LocalMux I__4424 (
            .O(N__27635),
            .I(N__27631));
    InMux I__4423 (
            .O(N__27634),
            .I(N__27628));
    Odrv4 I__4422 (
            .O(N__27631),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    LocalMux I__4421 (
            .O(N__27628),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    InMux I__4420 (
            .O(N__27623),
            .I(N__27619));
    InMux I__4419 (
            .O(N__27622),
            .I(N__27616));
    LocalMux I__4418 (
            .O(N__27619),
            .I(N__27613));
    LocalMux I__4417 (
            .O(N__27616),
            .I(N__27610));
    Span12Mux_v I__4416 (
            .O(N__27613),
            .I(N__27607));
    Span4Mux_v I__4415 (
            .O(N__27610),
            .I(N__27604));
    Odrv12 I__4414 (
            .O(N__27607),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    Odrv4 I__4413 (
            .O(N__27604),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    InMux I__4412 (
            .O(N__27599),
            .I(N__27595));
    CascadeMux I__4411 (
            .O(N__27598),
            .I(N__27591));
    LocalMux I__4410 (
            .O(N__27595),
            .I(N__27588));
    InMux I__4409 (
            .O(N__27594),
            .I(N__27585));
    InMux I__4408 (
            .O(N__27591),
            .I(N__27582));
    Span4Mux_h I__4407 (
            .O(N__27588),
            .I(N__27579));
    LocalMux I__4406 (
            .O(N__27585),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__4405 (
            .O(N__27582),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__4404 (
            .O(N__27579),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    CascadeMux I__4403 (
            .O(N__27572),
            .I(N__27569));
    InMux I__4402 (
            .O(N__27569),
            .I(N__27566));
    LocalMux I__4401 (
            .O(N__27566),
            .I(N__27561));
    InMux I__4400 (
            .O(N__27565),
            .I(N__27558));
    InMux I__4399 (
            .O(N__27564),
            .I(N__27555));
    Span4Mux_h I__4398 (
            .O(N__27561),
            .I(N__27552));
    LocalMux I__4397 (
            .O(N__27558),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__4396 (
            .O(N__27555),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__4395 (
            .O(N__27552),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__4394 (
            .O(N__27545),
            .I(N__27541));
    InMux I__4393 (
            .O(N__27544),
            .I(N__27538));
    LocalMux I__4392 (
            .O(N__27541),
            .I(N__27535));
    LocalMux I__4391 (
            .O(N__27538),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    Odrv4 I__4390 (
            .O(N__27535),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    InMux I__4389 (
            .O(N__27530),
            .I(N__27527));
    LocalMux I__4388 (
            .O(N__27527),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    InMux I__4387 (
            .O(N__27524),
            .I(N__27521));
    LocalMux I__4386 (
            .O(N__27521),
            .I(N__27516));
    InMux I__4385 (
            .O(N__27520),
            .I(N__27513));
    InMux I__4384 (
            .O(N__27519),
            .I(N__27510));
    Span4Mux_h I__4383 (
            .O(N__27516),
            .I(N__27505));
    LocalMux I__4382 (
            .O(N__27513),
            .I(N__27505));
    LocalMux I__4381 (
            .O(N__27510),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__4380 (
            .O(N__27505),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    CascadeMux I__4379 (
            .O(N__27500),
            .I(N__27497));
    InMux I__4378 (
            .O(N__27497),
            .I(N__27493));
    CascadeMux I__4377 (
            .O(N__27496),
            .I(N__27490));
    LocalMux I__4376 (
            .O(N__27493),
            .I(N__27486));
    InMux I__4375 (
            .O(N__27490),
            .I(N__27483));
    InMux I__4374 (
            .O(N__27489),
            .I(N__27480));
    Span4Mux_h I__4373 (
            .O(N__27486),
            .I(N__27475));
    LocalMux I__4372 (
            .O(N__27483),
            .I(N__27475));
    LocalMux I__4371 (
            .O(N__27480),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__4370 (
            .O(N__27475),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__4369 (
            .O(N__27470),
            .I(N__27467));
    LocalMux I__4368 (
            .O(N__27467),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    InMux I__4367 (
            .O(N__27464),
            .I(N__27460));
    InMux I__4366 (
            .O(N__27463),
            .I(N__27457));
    LocalMux I__4365 (
            .O(N__27460),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    LocalMux I__4364 (
            .O(N__27457),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    InMux I__4363 (
            .O(N__27452),
            .I(N__27446));
    InMux I__4362 (
            .O(N__27451),
            .I(N__27446));
    LocalMux I__4361 (
            .O(N__27446),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__4360 (
            .O(N__27443),
            .I(N__27440));
    InMux I__4359 (
            .O(N__27440),
            .I(N__27434));
    InMux I__4358 (
            .O(N__27439),
            .I(N__27434));
    LocalMux I__4357 (
            .O(N__27434),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__4356 (
            .O(N__27431),
            .I(N__27428));
    InMux I__4355 (
            .O(N__27428),
            .I(N__27425));
    LocalMux I__4354 (
            .O(N__27425),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    InMux I__4353 (
            .O(N__27422),
            .I(N__27419));
    LocalMux I__4352 (
            .O(N__27419),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    InMux I__4351 (
            .O(N__27416),
            .I(N__27412));
    InMux I__4350 (
            .O(N__27415),
            .I(N__27409));
    LocalMux I__4349 (
            .O(N__27412),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    LocalMux I__4348 (
            .O(N__27409),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    CascadeMux I__4347 (
            .O(N__27404),
            .I(N__27401));
    InMux I__4346 (
            .O(N__27401),
            .I(N__27398));
    LocalMux I__4345 (
            .O(N__27398),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    InMux I__4344 (
            .O(N__27395),
            .I(N__27391));
    InMux I__4343 (
            .O(N__27394),
            .I(N__27387));
    LocalMux I__4342 (
            .O(N__27391),
            .I(N__27384));
    InMux I__4341 (
            .O(N__27390),
            .I(N__27381));
    LocalMux I__4340 (
            .O(N__27387),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__4339 (
            .O(N__27384),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__4338 (
            .O(N__27381),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__4337 (
            .O(N__27374),
            .I(N__27371));
    LocalMux I__4336 (
            .O(N__27371),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__4335 (
            .O(N__27368),
            .I(N__27365));
    InMux I__4334 (
            .O(N__27365),
            .I(N__27362));
    LocalMux I__4333 (
            .O(N__27362),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__4332 (
            .O(N__27359),
            .I(N__27353));
    InMux I__4331 (
            .O(N__27358),
            .I(N__27353));
    LocalMux I__4330 (
            .O(N__27353),
            .I(N__27350));
    Odrv12 I__4329 (
            .O(N__27350),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    InMux I__4328 (
            .O(N__27347),
            .I(N__27343));
    InMux I__4327 (
            .O(N__27346),
            .I(N__27340));
    LocalMux I__4326 (
            .O(N__27343),
            .I(N__27335));
    LocalMux I__4325 (
            .O(N__27340),
            .I(N__27335));
    Odrv4 I__4324 (
            .O(N__27335),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    CascadeMux I__4323 (
            .O(N__27332),
            .I(N__27329));
    InMux I__4322 (
            .O(N__27329),
            .I(N__27325));
    InMux I__4321 (
            .O(N__27328),
            .I(N__27322));
    LocalMux I__4320 (
            .O(N__27325),
            .I(N__27316));
    LocalMux I__4319 (
            .O(N__27322),
            .I(N__27316));
    InMux I__4318 (
            .O(N__27321),
            .I(N__27313));
    Span4Mux_h I__4317 (
            .O(N__27316),
            .I(N__27310));
    LocalMux I__4316 (
            .O(N__27313),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__4315 (
            .O(N__27310),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    CascadeMux I__4314 (
            .O(N__27305),
            .I(N__27301));
    InMux I__4313 (
            .O(N__27304),
            .I(N__27296));
    InMux I__4312 (
            .O(N__27301),
            .I(N__27296));
    LocalMux I__4311 (
            .O(N__27296),
            .I(N__27292));
    InMux I__4310 (
            .O(N__27295),
            .I(N__27289));
    Span4Mux_h I__4309 (
            .O(N__27292),
            .I(N__27286));
    LocalMux I__4308 (
            .O(N__27289),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__4307 (
            .O(N__27286),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__4306 (
            .O(N__27281),
            .I(N__27278));
    LocalMux I__4305 (
            .O(N__27278),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    InMux I__4304 (
            .O(N__27275),
            .I(N__27271));
    InMux I__4303 (
            .O(N__27274),
            .I(N__27267));
    LocalMux I__4302 (
            .O(N__27271),
            .I(N__27264));
    InMux I__4301 (
            .O(N__27270),
            .I(N__27261));
    LocalMux I__4300 (
            .O(N__27267),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    Odrv12 I__4299 (
            .O(N__27264),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    LocalMux I__4298 (
            .O(N__27261),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    CascadeMux I__4297 (
            .O(N__27254),
            .I(elapsed_time_ns_1_RNI2COBB_0_15_cascade_));
    InMux I__4296 (
            .O(N__27251),
            .I(N__27248));
    LocalMux I__4295 (
            .O(N__27248),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    InMux I__4294 (
            .O(N__27245),
            .I(N__27239));
    InMux I__4293 (
            .O(N__27244),
            .I(N__27239));
    LocalMux I__4292 (
            .O(N__27239),
            .I(N__27235));
    InMux I__4291 (
            .O(N__27238),
            .I(N__27232));
    Span4Mux_h I__4290 (
            .O(N__27235),
            .I(N__27229));
    LocalMux I__4289 (
            .O(N__27232),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__4288 (
            .O(N__27229),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__4287 (
            .O(N__27224),
            .I(N__27221));
    InMux I__4286 (
            .O(N__27221),
            .I(N__27215));
    InMux I__4285 (
            .O(N__27220),
            .I(N__27215));
    LocalMux I__4284 (
            .O(N__27215),
            .I(N__27212));
    Span4Mux_h I__4283 (
            .O(N__27212),
            .I(N__27208));
    InMux I__4282 (
            .O(N__27211),
            .I(N__27205));
    Span4Mux_h I__4281 (
            .O(N__27208),
            .I(N__27202));
    LocalMux I__4280 (
            .O(N__27205),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__4279 (
            .O(N__27202),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__4278 (
            .O(N__27197),
            .I(N__27194));
    InMux I__4277 (
            .O(N__27194),
            .I(N__27191));
    LocalMux I__4276 (
            .O(N__27191),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    InMux I__4275 (
            .O(N__27188),
            .I(N__27184));
    InMux I__4274 (
            .O(N__27187),
            .I(N__27181));
    LocalMux I__4273 (
            .O(N__27184),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__4272 (
            .O(N__27181),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    CascadeMux I__4271 (
            .O(N__27176),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_));
    InMux I__4270 (
            .O(N__27173),
            .I(N__27169));
    InMux I__4269 (
            .O(N__27172),
            .I(N__27166));
    LocalMux I__4268 (
            .O(N__27169),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    LocalMux I__4267 (
            .O(N__27166),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    CascadeMux I__4266 (
            .O(N__27161),
            .I(elapsed_time_ns_1_RNILK91B_0_9_cascade_));
    InMux I__4265 (
            .O(N__27158),
            .I(N__27155));
    LocalMux I__4264 (
            .O(N__27155),
            .I(N__27152));
    Span4Mux_h I__4263 (
            .O(N__27152),
            .I(N__27149));
    Odrv4 I__4262 (
            .O(N__27149),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    InMux I__4261 (
            .O(N__27146),
            .I(N__27143));
    LocalMux I__4260 (
            .O(N__27143),
            .I(N__27140));
    Span4Mux_v I__4259 (
            .O(N__27140),
            .I(N__27137));
    Span4Mux_h I__4258 (
            .O(N__27137),
            .I(N__27134));
    Sp12to4 I__4257 (
            .O(N__27134),
            .I(N__27131));
    Span12Mux_h I__4256 (
            .O(N__27131),
            .I(N__27128));
    Odrv12 I__4255 (
            .O(N__27128),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__4254 (
            .O(N__27125),
            .I(N__27122));
    LocalMux I__4253 (
            .O(N__27122),
            .I(N__27117));
    CascadeMux I__4252 (
            .O(N__27121),
            .I(N__27107));
    CascadeMux I__4251 (
            .O(N__27120),
            .I(N__27104));
    Span4Mux_v I__4250 (
            .O(N__27117),
            .I(N__27101));
    CascadeMux I__4249 (
            .O(N__27116),
            .I(N__27098));
    CascadeMux I__4248 (
            .O(N__27115),
            .I(N__27095));
    CascadeMux I__4247 (
            .O(N__27114),
            .I(N__27091));
    CascadeMux I__4246 (
            .O(N__27113),
            .I(N__27087));
    CascadeMux I__4245 (
            .O(N__27112),
            .I(N__27084));
    CascadeMux I__4244 (
            .O(N__27111),
            .I(N__27081));
    CascadeMux I__4243 (
            .O(N__27110),
            .I(N__27078));
    InMux I__4242 (
            .O(N__27107),
            .I(N__27073));
    InMux I__4241 (
            .O(N__27104),
            .I(N__27073));
    Span4Mux_h I__4240 (
            .O(N__27101),
            .I(N__27070));
    InMux I__4239 (
            .O(N__27098),
            .I(N__27059));
    InMux I__4238 (
            .O(N__27095),
            .I(N__27059));
    InMux I__4237 (
            .O(N__27094),
            .I(N__27059));
    InMux I__4236 (
            .O(N__27091),
            .I(N__27059));
    InMux I__4235 (
            .O(N__27090),
            .I(N__27059));
    InMux I__4234 (
            .O(N__27087),
            .I(N__27054));
    InMux I__4233 (
            .O(N__27084),
            .I(N__27054));
    InMux I__4232 (
            .O(N__27081),
            .I(N__27049));
    InMux I__4231 (
            .O(N__27078),
            .I(N__27049));
    LocalMux I__4230 (
            .O(N__27073),
            .I(N__27038));
    Sp12to4 I__4229 (
            .O(N__27070),
            .I(N__27038));
    LocalMux I__4228 (
            .O(N__27059),
            .I(N__27038));
    LocalMux I__4227 (
            .O(N__27054),
            .I(N__27038));
    LocalMux I__4226 (
            .O(N__27049),
            .I(N__27038));
    Span12Mux_v I__4225 (
            .O(N__27038),
            .I(N__27035));
    Odrv12 I__4224 (
            .O(N__27035),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    InMux I__4223 (
            .O(N__27032),
            .I(N__27029));
    LocalMux I__4222 (
            .O(N__27029),
            .I(N__27026));
    Span4Mux_h I__4221 (
            .O(N__27026),
            .I(N__27023));
    Odrv4 I__4220 (
            .O(N__27023),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    InMux I__4219 (
            .O(N__27020),
            .I(N__27017));
    LocalMux I__4218 (
            .O(N__27017),
            .I(N__27014));
    Odrv4 I__4217 (
            .O(N__27014),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    InMux I__4216 (
            .O(N__27011),
            .I(N__27008));
    LocalMux I__4215 (
            .O(N__27008),
            .I(N__27005));
    Odrv12 I__4214 (
            .O(N__27005),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    InMux I__4213 (
            .O(N__27002),
            .I(N__26999));
    LocalMux I__4212 (
            .O(N__26999),
            .I(N__26996));
    Odrv4 I__4211 (
            .O(N__26996),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    InMux I__4210 (
            .O(N__26993),
            .I(N__26990));
    LocalMux I__4209 (
            .O(N__26990),
            .I(N__26987));
    Odrv4 I__4208 (
            .O(N__26987),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    InMux I__4207 (
            .O(N__26984),
            .I(N__26981));
    LocalMux I__4206 (
            .O(N__26981),
            .I(N__26978));
    Odrv12 I__4205 (
            .O(N__26978),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ));
    CascadeMux I__4204 (
            .O(N__26975),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8_cascade_));
    CascadeMux I__4203 (
            .O(N__26972),
            .I(N__26969));
    InMux I__4202 (
            .O(N__26969),
            .I(N__26966));
    LocalMux I__4201 (
            .O(N__26966),
            .I(N__26963));
    Odrv12 I__4200 (
            .O(N__26963),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__4199 (
            .O(N__26960),
            .I(N__26957));
    InMux I__4198 (
            .O(N__26957),
            .I(N__26954));
    LocalMux I__4197 (
            .O(N__26954),
            .I(N__26951));
    Odrv4 I__4196 (
            .O(N__26951),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    CascadeMux I__4195 (
            .O(N__26948),
            .I(N__26943));
    InMux I__4194 (
            .O(N__26947),
            .I(N__26940));
    InMux I__4193 (
            .O(N__26946),
            .I(N__26935));
    InMux I__4192 (
            .O(N__26943),
            .I(N__26935));
    LocalMux I__4191 (
            .O(N__26940),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__4190 (
            .O(N__26935),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__4189 (
            .O(N__26930),
            .I(N__26925));
    InMux I__4188 (
            .O(N__26929),
            .I(N__26920));
    InMux I__4187 (
            .O(N__26928),
            .I(N__26920));
    LocalMux I__4186 (
            .O(N__26925),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__4185 (
            .O(N__26920),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__4184 (
            .O(N__26915),
            .I(N__26912));
    LocalMux I__4183 (
            .O(N__26912),
            .I(N__26909));
    Odrv4 I__4182 (
            .O(N__26909),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    InMux I__4181 (
            .O(N__26906),
            .I(N__26900));
    InMux I__4180 (
            .O(N__26905),
            .I(N__26900));
    LocalMux I__4179 (
            .O(N__26900),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    CascadeMux I__4178 (
            .O(N__26897),
            .I(N__26893));
    InMux I__4177 (
            .O(N__26896),
            .I(N__26888));
    InMux I__4176 (
            .O(N__26893),
            .I(N__26888));
    LocalMux I__4175 (
            .O(N__26888),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    CascadeMux I__4174 (
            .O(N__26885),
            .I(N__26882));
    InMux I__4173 (
            .O(N__26882),
            .I(N__26879));
    LocalMux I__4172 (
            .O(N__26879),
            .I(N__26876));
    Span4Mux_h I__4171 (
            .O(N__26876),
            .I(N__26873));
    Odrv4 I__4170 (
            .O(N__26873),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    CascadeMux I__4169 (
            .O(N__26870),
            .I(N__26867));
    InMux I__4168 (
            .O(N__26867),
            .I(N__26864));
    LocalMux I__4167 (
            .O(N__26864),
            .I(N__26861));
    Span4Mux_v I__4166 (
            .O(N__26861),
            .I(N__26858));
    Odrv4 I__4165 (
            .O(N__26858),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    InMux I__4164 (
            .O(N__26855),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    InMux I__4163 (
            .O(N__26852),
            .I(N__26849));
    LocalMux I__4162 (
            .O(N__26849),
            .I(N__26846));
    Odrv4 I__4161 (
            .O(N__26846),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    CascadeMux I__4160 (
            .O(N__26843),
            .I(N__26838));
    InMux I__4159 (
            .O(N__26842),
            .I(N__26835));
    InMux I__4158 (
            .O(N__26841),
            .I(N__26830));
    InMux I__4157 (
            .O(N__26838),
            .I(N__26830));
    LocalMux I__4156 (
            .O(N__26835),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    LocalMux I__4155 (
            .O(N__26830),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    CascadeMux I__4154 (
            .O(N__26825),
            .I(N__26820));
    InMux I__4153 (
            .O(N__26824),
            .I(N__26817));
    InMux I__4152 (
            .O(N__26823),
            .I(N__26812));
    InMux I__4151 (
            .O(N__26820),
            .I(N__26812));
    LocalMux I__4150 (
            .O(N__26817),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    LocalMux I__4149 (
            .O(N__26812),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    CascadeMux I__4148 (
            .O(N__26807),
            .I(N__26804));
    InMux I__4147 (
            .O(N__26804),
            .I(N__26801));
    LocalMux I__4146 (
            .O(N__26801),
            .I(N__26798));
    Odrv4 I__4145 (
            .O(N__26798),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    InMux I__4144 (
            .O(N__26795),
            .I(N__26789));
    InMux I__4143 (
            .O(N__26794),
            .I(N__26789));
    LocalMux I__4142 (
            .O(N__26789),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    InMux I__4141 (
            .O(N__26786),
            .I(N__26780));
    InMux I__4140 (
            .O(N__26785),
            .I(N__26780));
    LocalMux I__4139 (
            .O(N__26780),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    InMux I__4138 (
            .O(N__26777),
            .I(N__26774));
    LocalMux I__4137 (
            .O(N__26774),
            .I(N__26771));
    Odrv4 I__4136 (
            .O(N__26771),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    InMux I__4135 (
            .O(N__26768),
            .I(N__26764));
    InMux I__4134 (
            .O(N__26767),
            .I(N__26761));
    LocalMux I__4133 (
            .O(N__26764),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__4132 (
            .O(N__26761),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__4131 (
            .O(N__26756),
            .I(N__26753));
    LocalMux I__4130 (
            .O(N__26753),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__4129 (
            .O(N__26750),
            .I(N__26746));
    InMux I__4128 (
            .O(N__26749),
            .I(N__26743));
    LocalMux I__4127 (
            .O(N__26746),
            .I(N__26740));
    LocalMux I__4126 (
            .O(N__26743),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__4125 (
            .O(N__26740),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__4124 (
            .O(N__26735),
            .I(N__26732));
    InMux I__4123 (
            .O(N__26732),
            .I(N__26729));
    LocalMux I__4122 (
            .O(N__26729),
            .I(N__26726));
    Odrv4 I__4121 (
            .O(N__26726),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__4120 (
            .O(N__26723),
            .I(N__26719));
    InMux I__4119 (
            .O(N__26722),
            .I(N__26716));
    LocalMux I__4118 (
            .O(N__26719),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__4117 (
            .O(N__26716),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__4116 (
            .O(N__26711),
            .I(N__26708));
    LocalMux I__4115 (
            .O(N__26708),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__4114 (
            .O(N__26705),
            .I(N__26702));
    LocalMux I__4113 (
            .O(N__26702),
            .I(N__26699));
    Span4Mux_v I__4112 (
            .O(N__26699),
            .I(N__26696));
    Odrv4 I__4111 (
            .O(N__26696),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    CascadeMux I__4110 (
            .O(N__26693),
            .I(N__26690));
    InMux I__4109 (
            .O(N__26690),
            .I(N__26687));
    LocalMux I__4108 (
            .O(N__26687),
            .I(N__26684));
    Span4Mux_v I__4107 (
            .O(N__26684),
            .I(N__26681));
    Odrv4 I__4106 (
            .O(N__26681),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    InMux I__4105 (
            .O(N__26678),
            .I(N__26675));
    LocalMux I__4104 (
            .O(N__26675),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    InMux I__4103 (
            .O(N__26672),
            .I(N__26668));
    InMux I__4102 (
            .O(N__26671),
            .I(N__26665));
    LocalMux I__4101 (
            .O(N__26668),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__4100 (
            .O(N__26665),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__4099 (
            .O(N__26660),
            .I(N__26657));
    InMux I__4098 (
            .O(N__26657),
            .I(N__26654));
    LocalMux I__4097 (
            .O(N__26654),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__4096 (
            .O(N__26651),
            .I(N__26647));
    InMux I__4095 (
            .O(N__26650),
            .I(N__26644));
    LocalMux I__4094 (
            .O(N__26647),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__4093 (
            .O(N__26644),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__4092 (
            .O(N__26639),
            .I(N__26636));
    InMux I__4091 (
            .O(N__26636),
            .I(N__26633));
    LocalMux I__4090 (
            .O(N__26633),
            .I(N__26630));
    Odrv4 I__4089 (
            .O(N__26630),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__4088 (
            .O(N__26627),
            .I(N__26624));
    LocalMux I__4087 (
            .O(N__26624),
            .I(N__26621));
    Odrv4 I__4086 (
            .O(N__26621),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__4085 (
            .O(N__26618),
            .I(N__26614));
    InMux I__4084 (
            .O(N__26617),
            .I(N__26611));
    LocalMux I__4083 (
            .O(N__26614),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__4082 (
            .O(N__26611),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__4081 (
            .O(N__26606),
            .I(N__26603));
    InMux I__4080 (
            .O(N__26603),
            .I(N__26600));
    LocalMux I__4079 (
            .O(N__26600),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    InMux I__4078 (
            .O(N__26597),
            .I(N__26593));
    InMux I__4077 (
            .O(N__26596),
            .I(N__26590));
    LocalMux I__4076 (
            .O(N__26593),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__4075 (
            .O(N__26590),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__4074 (
            .O(N__26585),
            .I(N__26582));
    LocalMux I__4073 (
            .O(N__26582),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__4072 (
            .O(N__26579),
            .I(N__26576));
    LocalMux I__4071 (
            .O(N__26576),
            .I(N__26573));
    Odrv4 I__4070 (
            .O(N__26573),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    InMux I__4069 (
            .O(N__26570),
            .I(N__26566));
    InMux I__4068 (
            .O(N__26569),
            .I(N__26563));
    LocalMux I__4067 (
            .O(N__26566),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__4066 (
            .O(N__26563),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__4065 (
            .O(N__26558),
            .I(N__26555));
    InMux I__4064 (
            .O(N__26555),
            .I(N__26552));
    LocalMux I__4063 (
            .O(N__26552),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__4062 (
            .O(N__26549),
            .I(N__26546));
    InMux I__4061 (
            .O(N__26546),
            .I(N__26543));
    LocalMux I__4060 (
            .O(N__26543),
            .I(N__26540));
    Odrv12 I__4059 (
            .O(N__26540),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    InMux I__4058 (
            .O(N__26537),
            .I(N__26533));
    InMux I__4057 (
            .O(N__26536),
            .I(N__26530));
    LocalMux I__4056 (
            .O(N__26533),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__4055 (
            .O(N__26530),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__4054 (
            .O(N__26525),
            .I(N__26522));
    LocalMux I__4053 (
            .O(N__26522),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__4052 (
            .O(N__26519),
            .I(N__26515));
    InMux I__4051 (
            .O(N__26518),
            .I(N__26512));
    LocalMux I__4050 (
            .O(N__26515),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__4049 (
            .O(N__26512),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__4048 (
            .O(N__26507),
            .I(N__26504));
    LocalMux I__4047 (
            .O(N__26504),
            .I(N__26501));
    Odrv12 I__4046 (
            .O(N__26501),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__4045 (
            .O(N__26498),
            .I(N__26495));
    InMux I__4044 (
            .O(N__26495),
            .I(N__26492));
    LocalMux I__4043 (
            .O(N__26492),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__4042 (
            .O(N__26489),
            .I(N__26485));
    InMux I__4041 (
            .O(N__26488),
            .I(N__26482));
    LocalMux I__4040 (
            .O(N__26485),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__4039 (
            .O(N__26482),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__4038 (
            .O(N__26477),
            .I(N__26474));
    InMux I__4037 (
            .O(N__26474),
            .I(N__26471));
    LocalMux I__4036 (
            .O(N__26471),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__4035 (
            .O(N__26468),
            .I(N__26465));
    InMux I__4034 (
            .O(N__26465),
            .I(N__26459));
    InMux I__4033 (
            .O(N__26464),
            .I(N__26459));
    LocalMux I__4032 (
            .O(N__26459),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__4031 (
            .O(N__26456),
            .I(N__26452));
    InMux I__4030 (
            .O(N__26455),
            .I(N__26449));
    LocalMux I__4029 (
            .O(N__26452),
            .I(N__26444));
    LocalMux I__4028 (
            .O(N__26449),
            .I(N__26444));
    Span4Mux_h I__4027 (
            .O(N__26444),
            .I(N__26440));
    CascadeMux I__4026 (
            .O(N__26443),
            .I(N__26437));
    Span4Mux_v I__4025 (
            .O(N__26440),
            .I(N__26434));
    InMux I__4024 (
            .O(N__26437),
            .I(N__26431));
    Span4Mux_v I__4023 (
            .O(N__26434),
            .I(N__26428));
    LocalMux I__4022 (
            .O(N__26431),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__4021 (
            .O(N__26428),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__4020 (
            .O(N__26423),
            .I(N__26420));
    InMux I__4019 (
            .O(N__26420),
            .I(N__26417));
    LocalMux I__4018 (
            .O(N__26417),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__4017 (
            .O(N__26414),
            .I(N__26410));
    InMux I__4016 (
            .O(N__26413),
            .I(N__26407));
    LocalMux I__4015 (
            .O(N__26410),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__4014 (
            .O(N__26407),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__4013 (
            .O(N__26402),
            .I(N__26399));
    LocalMux I__4012 (
            .O(N__26399),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__4011 (
            .O(N__26396),
            .I(N__26393));
    InMux I__4010 (
            .O(N__26393),
            .I(N__26390));
    LocalMux I__4009 (
            .O(N__26390),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__4008 (
            .O(N__26387),
            .I(N__26384));
    LocalMux I__4007 (
            .O(N__26384),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    InMux I__4006 (
            .O(N__26381),
            .I(N__26377));
    InMux I__4005 (
            .O(N__26380),
            .I(N__26374));
    LocalMux I__4004 (
            .O(N__26377),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__4003 (
            .O(N__26374),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__4002 (
            .O(N__26369),
            .I(N__26366));
    InMux I__4001 (
            .O(N__26366),
            .I(N__26363));
    LocalMux I__4000 (
            .O(N__26363),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__3999 (
            .O(N__26360),
            .I(N__26357));
    InMux I__3998 (
            .O(N__26357),
            .I(N__26354));
    LocalMux I__3997 (
            .O(N__26354),
            .I(N__26351));
    Odrv4 I__3996 (
            .O(N__26351),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    InMux I__3995 (
            .O(N__26348),
            .I(N__26344));
    InMux I__3994 (
            .O(N__26347),
            .I(N__26341));
    LocalMux I__3993 (
            .O(N__26344),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__3992 (
            .O(N__26341),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__3991 (
            .O(N__26336),
            .I(N__26333));
    LocalMux I__3990 (
            .O(N__26333),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__3989 (
            .O(N__26330),
            .I(N__26324));
    InMux I__3988 (
            .O(N__26329),
            .I(N__26324));
    LocalMux I__3987 (
            .O(N__26324),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    InMux I__3986 (
            .O(N__26321),
            .I(N__26314));
    InMux I__3985 (
            .O(N__26320),
            .I(N__26314));
    InMux I__3984 (
            .O(N__26319),
            .I(N__26311));
    LocalMux I__3983 (
            .O(N__26314),
            .I(N__26308));
    LocalMux I__3982 (
            .O(N__26311),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__3981 (
            .O(N__26308),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__3980 (
            .O(N__26303),
            .I(N__26300));
    InMux I__3979 (
            .O(N__26300),
            .I(N__26293));
    InMux I__3978 (
            .O(N__26299),
            .I(N__26293));
    InMux I__3977 (
            .O(N__26298),
            .I(N__26290));
    LocalMux I__3976 (
            .O(N__26293),
            .I(N__26287));
    LocalMux I__3975 (
            .O(N__26290),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__3974 (
            .O(N__26287),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__3973 (
            .O(N__26282),
            .I(N__26279));
    LocalMux I__3972 (
            .O(N__26279),
            .I(N__26276));
    Odrv4 I__3971 (
            .O(N__26276),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__3970 (
            .O(N__26273),
            .I(N__26270));
    LocalMux I__3969 (
            .O(N__26270),
            .I(N__26267));
    Odrv4 I__3968 (
            .O(N__26267),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__3967 (
            .O(N__26264),
            .I(N__26261));
    LocalMux I__3966 (
            .O(N__26261),
            .I(N__26258));
    Odrv4 I__3965 (
            .O(N__26258),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__3964 (
            .O(N__26255),
            .I(N__26252));
    LocalMux I__3963 (
            .O(N__26252),
            .I(N__26249));
    Odrv4 I__3962 (
            .O(N__26249),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    InMux I__3961 (
            .O(N__26246),
            .I(N__26243));
    LocalMux I__3960 (
            .O(N__26243),
            .I(N__26240));
    Odrv4 I__3959 (
            .O(N__26240),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    InMux I__3958 (
            .O(N__26237),
            .I(N__26234));
    LocalMux I__3957 (
            .O(N__26234),
            .I(N__26231));
    Odrv12 I__3956 (
            .O(N__26231),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    InMux I__3955 (
            .O(N__26228),
            .I(N__26225));
    LocalMux I__3954 (
            .O(N__26225),
            .I(N__26222));
    Span12Mux_v I__3953 (
            .O(N__26222),
            .I(N__26218));
    InMux I__3952 (
            .O(N__26221),
            .I(N__26215));
    Odrv12 I__3951 (
            .O(N__26218),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__3950 (
            .O(N__26215),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    IoInMux I__3949 (
            .O(N__26210),
            .I(N__26189));
    InMux I__3948 (
            .O(N__26209),
            .I(N__26182));
    InMux I__3947 (
            .O(N__26208),
            .I(N__26182));
    InMux I__3946 (
            .O(N__26207),
            .I(N__26182));
    InMux I__3945 (
            .O(N__26206),
            .I(N__26162));
    InMux I__3944 (
            .O(N__26205),
            .I(N__26162));
    InMux I__3943 (
            .O(N__26204),
            .I(N__26162));
    InMux I__3942 (
            .O(N__26203),
            .I(N__26153));
    InMux I__3941 (
            .O(N__26202),
            .I(N__26153));
    InMux I__3940 (
            .O(N__26201),
            .I(N__26153));
    InMux I__3939 (
            .O(N__26200),
            .I(N__26153));
    InMux I__3938 (
            .O(N__26199),
            .I(N__26144));
    InMux I__3937 (
            .O(N__26198),
            .I(N__26144));
    InMux I__3936 (
            .O(N__26197),
            .I(N__26144));
    InMux I__3935 (
            .O(N__26196),
            .I(N__26144));
    InMux I__3934 (
            .O(N__26195),
            .I(N__26135));
    InMux I__3933 (
            .O(N__26194),
            .I(N__26135));
    InMux I__3932 (
            .O(N__26193),
            .I(N__26135));
    InMux I__3931 (
            .O(N__26192),
            .I(N__26135));
    LocalMux I__3930 (
            .O(N__26189),
            .I(N__26132));
    LocalMux I__3929 (
            .O(N__26182),
            .I(N__26129));
    InMux I__3928 (
            .O(N__26181),
            .I(N__26126));
    InMux I__3927 (
            .O(N__26180),
            .I(N__26117));
    InMux I__3926 (
            .O(N__26179),
            .I(N__26117));
    InMux I__3925 (
            .O(N__26178),
            .I(N__26117));
    InMux I__3924 (
            .O(N__26177),
            .I(N__26117));
    InMux I__3923 (
            .O(N__26176),
            .I(N__26108));
    InMux I__3922 (
            .O(N__26175),
            .I(N__26108));
    InMux I__3921 (
            .O(N__26174),
            .I(N__26108));
    InMux I__3920 (
            .O(N__26173),
            .I(N__26108));
    InMux I__3919 (
            .O(N__26172),
            .I(N__26099));
    InMux I__3918 (
            .O(N__26171),
            .I(N__26099));
    InMux I__3917 (
            .O(N__26170),
            .I(N__26099));
    InMux I__3916 (
            .O(N__26169),
            .I(N__26099));
    LocalMux I__3915 (
            .O(N__26162),
            .I(N__26096));
    LocalMux I__3914 (
            .O(N__26153),
            .I(N__26091));
    LocalMux I__3913 (
            .O(N__26144),
            .I(N__26091));
    LocalMux I__3912 (
            .O(N__26135),
            .I(N__26088));
    Span12Mux_s2_v I__3911 (
            .O(N__26132),
            .I(N__26085));
    Span12Mux_v I__3910 (
            .O(N__26129),
            .I(N__26080));
    LocalMux I__3909 (
            .O(N__26126),
            .I(N__26080));
    LocalMux I__3908 (
            .O(N__26117),
            .I(N__26067));
    LocalMux I__3907 (
            .O(N__26108),
            .I(N__26067));
    LocalMux I__3906 (
            .O(N__26099),
            .I(N__26067));
    Span4Mux_v I__3905 (
            .O(N__26096),
            .I(N__26067));
    Span4Mux_v I__3904 (
            .O(N__26091),
            .I(N__26067));
    Span4Mux_h I__3903 (
            .O(N__26088),
            .I(N__26067));
    Span12Mux_v I__3902 (
            .O(N__26085),
            .I(N__26064));
    Odrv12 I__3901 (
            .O(N__26080),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__3900 (
            .O(N__26067),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv12 I__3899 (
            .O(N__26064),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__3898 (
            .O(N__26057),
            .I(N__26054));
    LocalMux I__3897 (
            .O(N__26054),
            .I(N__26051));
    Span4Mux_v I__3896 (
            .O(N__26051),
            .I(N__26048));
    Odrv4 I__3895 (
            .O(N__26048),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__3894 (
            .O(N__26045),
            .I(N__26042));
    LocalMux I__3893 (
            .O(N__26042),
            .I(N__26037));
    InMux I__3892 (
            .O(N__26041),
            .I(N__26032));
    InMux I__3891 (
            .O(N__26040),
            .I(N__26032));
    Odrv12 I__3890 (
            .O(N__26037),
            .I(\current_shift_inst.PI_CTRL.N_160 ));
    LocalMux I__3889 (
            .O(N__26032),
            .I(\current_shift_inst.PI_CTRL.N_160 ));
    InMux I__3888 (
            .O(N__26027),
            .I(N__26023));
    InMux I__3887 (
            .O(N__26026),
            .I(N__26020));
    LocalMux I__3886 (
            .O(N__26023),
            .I(N__26017));
    LocalMux I__3885 (
            .O(N__26020),
            .I(N__26014));
    Span4Mux_v I__3884 (
            .O(N__26017),
            .I(N__26009));
    Span4Mux_s3_h I__3883 (
            .O(N__26014),
            .I(N__26009));
    Span4Mux_h I__3882 (
            .O(N__26009),
            .I(N__26006));
    Odrv4 I__3881 (
            .O(N__26006),
            .I(pwm_duty_input_2));
    CascadeMux I__3880 (
            .O(N__26003),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__3879 (
            .O(N__26000),
            .I(N__25997));
    InMux I__3878 (
            .O(N__25997),
            .I(N__25992));
    CascadeMux I__3877 (
            .O(N__25996),
            .I(N__25989));
    InMux I__3876 (
            .O(N__25995),
            .I(N__25986));
    LocalMux I__3875 (
            .O(N__25992),
            .I(N__25982));
    InMux I__3874 (
            .O(N__25989),
            .I(N__25979));
    LocalMux I__3873 (
            .O(N__25986),
            .I(N__25976));
    InMux I__3872 (
            .O(N__25985),
            .I(N__25973));
    Odrv12 I__3871 (
            .O(N__25982),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__3870 (
            .O(N__25979),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__3869 (
            .O(N__25976),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__3868 (
            .O(N__25973),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    CascadeMux I__3867 (
            .O(N__25964),
            .I(N__25961));
    InMux I__3866 (
            .O(N__25961),
            .I(N__25958));
    LocalMux I__3865 (
            .O(N__25958),
            .I(N__25954));
    InMux I__3864 (
            .O(N__25957),
            .I(N__25950));
    Span4Mux_v I__3863 (
            .O(N__25954),
            .I(N__25946));
    InMux I__3862 (
            .O(N__25953),
            .I(N__25943));
    LocalMux I__3861 (
            .O(N__25950),
            .I(N__25940));
    InMux I__3860 (
            .O(N__25949),
            .I(N__25937));
    Odrv4 I__3859 (
            .O(N__25946),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__3858 (
            .O(N__25943),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__3857 (
            .O(N__25940),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__3856 (
            .O(N__25937),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    CascadeMux I__3855 (
            .O(N__25928),
            .I(N__25925));
    InMux I__3854 (
            .O(N__25925),
            .I(N__25921));
    CascadeMux I__3853 (
            .O(N__25924),
            .I(N__25918));
    LocalMux I__3852 (
            .O(N__25921),
            .I(N__25915));
    InMux I__3851 (
            .O(N__25918),
            .I(N__25911));
    Span4Mux_v I__3850 (
            .O(N__25915),
            .I(N__25907));
    InMux I__3849 (
            .O(N__25914),
            .I(N__25904));
    LocalMux I__3848 (
            .O(N__25911),
            .I(N__25901));
    InMux I__3847 (
            .O(N__25910),
            .I(N__25898));
    Odrv4 I__3846 (
            .O(N__25907),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__3845 (
            .O(N__25904),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv12 I__3844 (
            .O(N__25901),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__3843 (
            .O(N__25898),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    CascadeMux I__3842 (
            .O(N__25889),
            .I(N__25886));
    InMux I__3841 (
            .O(N__25886),
            .I(N__25883));
    LocalMux I__3840 (
            .O(N__25883),
            .I(N__25878));
    InMux I__3839 (
            .O(N__25882),
            .I(N__25874));
    CascadeMux I__3838 (
            .O(N__25881),
            .I(N__25871));
    Span4Mux_v I__3837 (
            .O(N__25878),
            .I(N__25868));
    InMux I__3836 (
            .O(N__25877),
            .I(N__25865));
    LocalMux I__3835 (
            .O(N__25874),
            .I(N__25862));
    InMux I__3834 (
            .O(N__25871),
            .I(N__25859));
    Odrv4 I__3833 (
            .O(N__25868),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__3832 (
            .O(N__25865),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__3831 (
            .O(N__25862),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__3830 (
            .O(N__25859),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    CascadeMux I__3829 (
            .O(N__25850),
            .I(N__25847));
    InMux I__3828 (
            .O(N__25847),
            .I(N__25844));
    LocalMux I__3827 (
            .O(N__25844),
            .I(N__25841));
    Span4Mux_h I__3826 (
            .O(N__25841),
            .I(N__25838));
    Odrv4 I__3825 (
            .O(N__25838),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__3824 (
            .O(N__25835),
            .I(N__25832));
    LocalMux I__3823 (
            .O(N__25832),
            .I(N__25829));
    Span12Mux_s7_h I__3822 (
            .O(N__25829),
            .I(N__25826));
    Odrv12 I__3821 (
            .O(N__25826),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__3820 (
            .O(N__25823),
            .I(N__25820));
    LocalMux I__3819 (
            .O(N__25820),
            .I(N__25817));
    Odrv4 I__3818 (
            .O(N__25817),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__3817 (
            .O(N__25814),
            .I(N__25811));
    LocalMux I__3816 (
            .O(N__25811),
            .I(N__25808));
    Span4Mux_h I__3815 (
            .O(N__25808),
            .I(N__25805));
    Odrv4 I__3814 (
            .O(N__25805),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__3813 (
            .O(N__25802),
            .I(N__25799));
    LocalMux I__3812 (
            .O(N__25799),
            .I(N__25796));
    Odrv12 I__3811 (
            .O(N__25796),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__3810 (
            .O(N__25793),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__3809 (
            .O(N__25790),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__3808 (
            .O(N__25787),
            .I(bfn_7_13_0_));
    InMux I__3807 (
            .O(N__25784),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__3806 (
            .O(N__25781),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__3805 (
            .O(N__25778),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__3804 (
            .O(N__25775),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__3803 (
            .O(N__25772),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__3802 (
            .O(N__25769),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__3801 (
            .O(N__25766),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__3800 (
            .O(N__25763),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__3799 (
            .O(N__25760),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__3798 (
            .O(N__25757),
            .I(bfn_7_12_0_));
    InMux I__3797 (
            .O(N__25754),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__3796 (
            .O(N__25751),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__3795 (
            .O(N__25748),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__3794 (
            .O(N__25745),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__3793 (
            .O(N__25742),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__3792 (
            .O(N__25739),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__3791 (
            .O(N__25736),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__3790 (
            .O(N__25733),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__3789 (
            .O(N__25730),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__3788 (
            .O(N__25727),
            .I(bfn_7_11_0_));
    InMux I__3787 (
            .O(N__25724),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__3786 (
            .O(N__25721),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__3785 (
            .O(N__25718),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__3784 (
            .O(N__25715),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    CascadeMux I__3783 (
            .O(N__25712),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ));
    InMux I__3782 (
            .O(N__25709),
            .I(N__25703));
    InMux I__3781 (
            .O(N__25708),
            .I(N__25703));
    LocalMux I__3780 (
            .O(N__25703),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    CascadeMux I__3779 (
            .O(N__25700),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__3778 (
            .O(N__25697),
            .I(N__25694));
    InMux I__3777 (
            .O(N__25694),
            .I(N__25691));
    LocalMux I__3776 (
            .O(N__25691),
            .I(N__25688));
    Odrv4 I__3775 (
            .O(N__25688),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__3774 (
            .O(N__25685),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__3773 (
            .O(N__25682),
            .I(N__25679));
    InMux I__3772 (
            .O(N__25679),
            .I(N__25676));
    LocalMux I__3771 (
            .O(N__25676),
            .I(N__25673));
    Odrv4 I__3770 (
            .O(N__25673),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ));
    InMux I__3769 (
            .O(N__25670),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__3768 (
            .O(N__25667),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__3767 (
            .O(N__25664),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__3766 (
            .O(N__25661),
            .I(N__25657));
    InMux I__3765 (
            .O(N__25660),
            .I(N__25654));
    LocalMux I__3764 (
            .O(N__25657),
            .I(N__25651));
    LocalMux I__3763 (
            .O(N__25654),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    Odrv4 I__3762 (
            .O(N__25651),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__3761 (
            .O(N__25646),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__3760 (
            .O(N__25643),
            .I(N__25640));
    LocalMux I__3759 (
            .O(N__25640),
            .I(N__25636));
    InMux I__3758 (
            .O(N__25639),
            .I(N__25633));
    Odrv4 I__3757 (
            .O(N__25636),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__3756 (
            .O(N__25633),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__3755 (
            .O(N__25628),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    CascadeMux I__3754 (
            .O(N__25625),
            .I(N__25622));
    InMux I__3753 (
            .O(N__25622),
            .I(N__25619));
    LocalMux I__3752 (
            .O(N__25619),
            .I(N__25613));
    InMux I__3751 (
            .O(N__25618),
            .I(N__25610));
    InMux I__3750 (
            .O(N__25617),
            .I(N__25607));
    InMux I__3749 (
            .O(N__25616),
            .I(N__25604));
    Span4Mux_v I__3748 (
            .O(N__25613),
            .I(N__25599));
    LocalMux I__3747 (
            .O(N__25610),
            .I(N__25599));
    LocalMux I__3746 (
            .O(N__25607),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__3745 (
            .O(N__25604),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__3744 (
            .O(N__25599),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__3743 (
            .O(N__25592),
            .I(N__25589));
    LocalMux I__3742 (
            .O(N__25589),
            .I(N__25585));
    InMux I__3741 (
            .O(N__25588),
            .I(N__25582));
    Odrv4 I__3740 (
            .O(N__25585),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__3739 (
            .O(N__25582),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__3738 (
            .O(N__25577),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__3737 (
            .O(N__25574),
            .I(N__25571));
    InMux I__3736 (
            .O(N__25571),
            .I(N__25568));
    LocalMux I__3735 (
            .O(N__25568),
            .I(N__25564));
    InMux I__3734 (
            .O(N__25567),
            .I(N__25560));
    Span4Mux_v I__3733 (
            .O(N__25564),
            .I(N__25556));
    InMux I__3732 (
            .O(N__25563),
            .I(N__25553));
    LocalMux I__3731 (
            .O(N__25560),
            .I(N__25550));
    InMux I__3730 (
            .O(N__25559),
            .I(N__25547));
    Odrv4 I__3729 (
            .O(N__25556),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__3728 (
            .O(N__25553),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__3727 (
            .O(N__25550),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__3726 (
            .O(N__25547),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__3725 (
            .O(N__25538),
            .I(N__25534));
    InMux I__3724 (
            .O(N__25537),
            .I(N__25531));
    LocalMux I__3723 (
            .O(N__25534),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    LocalMux I__3722 (
            .O(N__25531),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__3721 (
            .O(N__25526),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    CascadeMux I__3720 (
            .O(N__25523),
            .I(N__25518));
    InMux I__3719 (
            .O(N__25522),
            .I(N__25496));
    InMux I__3718 (
            .O(N__25521),
            .I(N__25496));
    InMux I__3717 (
            .O(N__25518),
            .I(N__25487));
    InMux I__3716 (
            .O(N__25517),
            .I(N__25487));
    InMux I__3715 (
            .O(N__25516),
            .I(N__25487));
    InMux I__3714 (
            .O(N__25515),
            .I(N__25487));
    InMux I__3713 (
            .O(N__25514),
            .I(N__25480));
    InMux I__3712 (
            .O(N__25513),
            .I(N__25480));
    InMux I__3711 (
            .O(N__25512),
            .I(N__25480));
    InMux I__3710 (
            .O(N__25511),
            .I(N__25476));
    InMux I__3709 (
            .O(N__25510),
            .I(N__25467));
    InMux I__3708 (
            .O(N__25509),
            .I(N__25462));
    InMux I__3707 (
            .O(N__25508),
            .I(N__25462));
    InMux I__3706 (
            .O(N__25507),
            .I(N__25447));
    InMux I__3705 (
            .O(N__25506),
            .I(N__25447));
    InMux I__3704 (
            .O(N__25505),
            .I(N__25447));
    InMux I__3703 (
            .O(N__25504),
            .I(N__25447));
    InMux I__3702 (
            .O(N__25503),
            .I(N__25447));
    InMux I__3701 (
            .O(N__25502),
            .I(N__25447));
    InMux I__3700 (
            .O(N__25501),
            .I(N__25447));
    LocalMux I__3699 (
            .O(N__25496),
            .I(N__25440));
    LocalMux I__3698 (
            .O(N__25487),
            .I(N__25440));
    LocalMux I__3697 (
            .O(N__25480),
            .I(N__25440));
    InMux I__3696 (
            .O(N__25479),
            .I(N__25437));
    LocalMux I__3695 (
            .O(N__25476),
            .I(N__25432));
    InMux I__3694 (
            .O(N__25475),
            .I(N__25419));
    InMux I__3693 (
            .O(N__25474),
            .I(N__25419));
    InMux I__3692 (
            .O(N__25473),
            .I(N__25419));
    InMux I__3691 (
            .O(N__25472),
            .I(N__25419));
    InMux I__3690 (
            .O(N__25471),
            .I(N__25419));
    InMux I__3689 (
            .O(N__25470),
            .I(N__25419));
    LocalMux I__3688 (
            .O(N__25467),
            .I(N__25414));
    LocalMux I__3687 (
            .O(N__25462),
            .I(N__25414));
    LocalMux I__3686 (
            .O(N__25447),
            .I(N__25409));
    Span4Mux_v I__3685 (
            .O(N__25440),
            .I(N__25409));
    LocalMux I__3684 (
            .O(N__25437),
            .I(N__25405));
    InMux I__3683 (
            .O(N__25436),
            .I(N__25398));
    InMux I__3682 (
            .O(N__25435),
            .I(N__25398));
    Span12Mux_s10_v I__3681 (
            .O(N__25432),
            .I(N__25393));
    LocalMux I__3680 (
            .O(N__25419),
            .I(N__25393));
    Span4Mux_v I__3679 (
            .O(N__25414),
            .I(N__25390));
    Sp12to4 I__3678 (
            .O(N__25409),
            .I(N__25387));
    InMux I__3677 (
            .O(N__25408),
            .I(N__25384));
    Span4Mux_h I__3676 (
            .O(N__25405),
            .I(N__25381));
    InMux I__3675 (
            .O(N__25404),
            .I(N__25378));
    InMux I__3674 (
            .O(N__25403),
            .I(N__25375));
    LocalMux I__3673 (
            .O(N__25398),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__3672 (
            .O(N__25393),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3671 (
            .O(N__25390),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__3670 (
            .O(N__25387),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3669 (
            .O(N__25384),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3668 (
            .O(N__25381),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3667 (
            .O(N__25378),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3666 (
            .O(N__25375),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__3665 (
            .O(N__25358),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    CascadeMux I__3664 (
            .O(N__25355),
            .I(N__25350));
    InMux I__3663 (
            .O(N__25354),
            .I(N__25347));
    InMux I__3662 (
            .O(N__25353),
            .I(N__25344));
    InMux I__3661 (
            .O(N__25350),
            .I(N__25341));
    LocalMux I__3660 (
            .O(N__25347),
            .I(N__25338));
    LocalMux I__3659 (
            .O(N__25344),
            .I(N__25335));
    LocalMux I__3658 (
            .O(N__25341),
            .I(N__25332));
    Span4Mux_h I__3657 (
            .O(N__25338),
            .I(N__25329));
    Span4Mux_h I__3656 (
            .O(N__25335),
            .I(N__25326));
    Odrv12 I__3655 (
            .O(N__25332),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__3654 (
            .O(N__25329),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__3653 (
            .O(N__25326),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__3652 (
            .O(N__25319),
            .I(N__25314));
    InMux I__3651 (
            .O(N__25318),
            .I(N__25309));
    InMux I__3650 (
            .O(N__25317),
            .I(N__25309));
    LocalMux I__3649 (
            .O(N__25314),
            .I(N__25306));
    LocalMux I__3648 (
            .O(N__25309),
            .I(N__25303));
    Span4Mux_s1_h I__3647 (
            .O(N__25306),
            .I(N__25300));
    Span4Mux_v I__3646 (
            .O(N__25303),
            .I(N__25297));
    Span4Mux_h I__3645 (
            .O(N__25300),
            .I(N__25294));
    Odrv4 I__3644 (
            .O(N__25297),
            .I(pwm_duty_input_8));
    Odrv4 I__3643 (
            .O(N__25294),
            .I(pwm_duty_input_8));
    InMux I__3642 (
            .O(N__25289),
            .I(N__25283));
    InMux I__3641 (
            .O(N__25288),
            .I(N__25283));
    LocalMux I__3640 (
            .O(N__25283),
            .I(N__25277));
    InMux I__3639 (
            .O(N__25282),
            .I(N__25270));
    InMux I__3638 (
            .O(N__25281),
            .I(N__25270));
    InMux I__3637 (
            .O(N__25280),
            .I(N__25270));
    Span4Mux_h I__3636 (
            .O(N__25277),
            .I(N__25263));
    LocalMux I__3635 (
            .O(N__25270),
            .I(N__25263));
    InMux I__3634 (
            .O(N__25269),
            .I(N__25260));
    InMux I__3633 (
            .O(N__25268),
            .I(N__25257));
    Odrv4 I__3632 (
            .O(N__25263),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    LocalMux I__3631 (
            .O(N__25260),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    LocalMux I__3630 (
            .O(N__25257),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    InMux I__3629 (
            .O(N__25250),
            .I(N__25247));
    LocalMux I__3628 (
            .O(N__25247),
            .I(N__25244));
    Span4Mux_v I__3627 (
            .O(N__25244),
            .I(N__25237));
    InMux I__3626 (
            .O(N__25243),
            .I(N__25228));
    InMux I__3625 (
            .O(N__25242),
            .I(N__25228));
    InMux I__3624 (
            .O(N__25241),
            .I(N__25228));
    CascadeMux I__3623 (
            .O(N__25240),
            .I(N__25224));
    Span4Mux_v I__3622 (
            .O(N__25237),
            .I(N__25221));
    InMux I__3621 (
            .O(N__25236),
            .I(N__25216));
    InMux I__3620 (
            .O(N__25235),
            .I(N__25216));
    LocalMux I__3619 (
            .O(N__25228),
            .I(N__25211));
    InMux I__3618 (
            .O(N__25227),
            .I(N__25206));
    InMux I__3617 (
            .O(N__25224),
            .I(N__25206));
    Span4Mux_v I__3616 (
            .O(N__25221),
            .I(N__25201));
    LocalMux I__3615 (
            .O(N__25216),
            .I(N__25201));
    InMux I__3614 (
            .O(N__25215),
            .I(N__25196));
    InMux I__3613 (
            .O(N__25214),
            .I(N__25196));
    Span4Mux_v I__3612 (
            .O(N__25211),
            .I(N__25191));
    LocalMux I__3611 (
            .O(N__25206),
            .I(N__25191));
    Span4Mux_h I__3610 (
            .O(N__25201),
            .I(N__25188));
    LocalMux I__3609 (
            .O(N__25196),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__3608 (
            .O(N__25191),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__3607 (
            .O(N__25188),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__3606 (
            .O(N__25181),
            .I(N__25176));
    InMux I__3605 (
            .O(N__25180),
            .I(N__25171));
    InMux I__3604 (
            .O(N__25179),
            .I(N__25171));
    InMux I__3603 (
            .O(N__25176),
            .I(N__25168));
    LocalMux I__3602 (
            .O(N__25171),
            .I(N__25165));
    LocalMux I__3601 (
            .O(N__25168),
            .I(N__25162));
    Span4Mux_h I__3600 (
            .O(N__25165),
            .I(N__25159));
    Odrv12 I__3599 (
            .O(N__25162),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__3598 (
            .O(N__25159),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    CascadeMux I__3597 (
            .O(N__25154),
            .I(N__25148));
    CascadeMux I__3596 (
            .O(N__25153),
            .I(N__25144));
    CascadeMux I__3595 (
            .O(N__25152),
            .I(N__25141));
    InMux I__3594 (
            .O(N__25151),
            .I(N__25136));
    InMux I__3593 (
            .O(N__25148),
            .I(N__25133));
    InMux I__3592 (
            .O(N__25147),
            .I(N__25126));
    InMux I__3591 (
            .O(N__25144),
            .I(N__25126));
    InMux I__3590 (
            .O(N__25141),
            .I(N__25126));
    InMux I__3589 (
            .O(N__25140),
            .I(N__25123));
    InMux I__3588 (
            .O(N__25139),
            .I(N__25120));
    LocalMux I__3587 (
            .O(N__25136),
            .I(\current_shift_inst.PI_CTRL.N_158 ));
    LocalMux I__3586 (
            .O(N__25133),
            .I(\current_shift_inst.PI_CTRL.N_158 ));
    LocalMux I__3585 (
            .O(N__25126),
            .I(\current_shift_inst.PI_CTRL.N_158 ));
    LocalMux I__3584 (
            .O(N__25123),
            .I(\current_shift_inst.PI_CTRL.N_158 ));
    LocalMux I__3583 (
            .O(N__25120),
            .I(\current_shift_inst.PI_CTRL.N_158 ));
    InMux I__3582 (
            .O(N__25109),
            .I(N__25102));
    InMux I__3581 (
            .O(N__25108),
            .I(N__25102));
    InMux I__3580 (
            .O(N__25107),
            .I(N__25099));
    LocalMux I__3579 (
            .O(N__25102),
            .I(N__25096));
    LocalMux I__3578 (
            .O(N__25099),
            .I(N__25093));
    Span4Mux_v I__3577 (
            .O(N__25096),
            .I(N__25090));
    Span12Mux_s7_v I__3576 (
            .O(N__25093),
            .I(N__25087));
    Odrv4 I__3575 (
            .O(N__25090),
            .I(pwm_duty_input_9));
    Odrv12 I__3574 (
            .O(N__25087),
            .I(pwm_duty_input_9));
    InMux I__3573 (
            .O(N__25082),
            .I(N__25079));
    LocalMux I__3572 (
            .O(N__25079),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    CascadeMux I__3571 (
            .O(N__25076),
            .I(N__25073));
    InMux I__3570 (
            .O(N__25073),
            .I(N__25070));
    LocalMux I__3569 (
            .O(N__25070),
            .I(N__25066));
    CascadeMux I__3568 (
            .O(N__25069),
            .I(N__25061));
    Span4Mux_v I__3567 (
            .O(N__25066),
            .I(N__25058));
    CascadeMux I__3566 (
            .O(N__25065),
            .I(N__25055));
    InMux I__3565 (
            .O(N__25064),
            .I(N__25052));
    InMux I__3564 (
            .O(N__25061),
            .I(N__25049));
    Span4Mux_v I__3563 (
            .O(N__25058),
            .I(N__25046));
    InMux I__3562 (
            .O(N__25055),
            .I(N__25043));
    LocalMux I__3561 (
            .O(N__25052),
            .I(N__25038));
    LocalMux I__3560 (
            .O(N__25049),
            .I(N__25038));
    Odrv4 I__3559 (
            .O(N__25046),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__3558 (
            .O(N__25043),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__3557 (
            .O(N__25038),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__3556 (
            .O(N__25031),
            .I(N__25025));
    InMux I__3555 (
            .O(N__25030),
            .I(N__25025));
    LocalMux I__3554 (
            .O(N__25025),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__3553 (
            .O(N__25022),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    CascadeMux I__3552 (
            .O(N__25019),
            .I(N__25016));
    InMux I__3551 (
            .O(N__25016),
            .I(N__25013));
    LocalMux I__3550 (
            .O(N__25013),
            .I(N__25007));
    InMux I__3549 (
            .O(N__25012),
            .I(N__25002));
    InMux I__3548 (
            .O(N__25011),
            .I(N__25002));
    InMux I__3547 (
            .O(N__25010),
            .I(N__24999));
    Span12Mux_v I__3546 (
            .O(N__25007),
            .I(N__24994));
    LocalMux I__3545 (
            .O(N__25002),
            .I(N__24994));
    LocalMux I__3544 (
            .O(N__24999),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv12 I__3543 (
            .O(N__24994),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__3542 (
            .O(N__24989),
            .I(N__24986));
    InMux I__3541 (
            .O(N__24986),
            .I(N__24980));
    InMux I__3540 (
            .O(N__24985),
            .I(N__24980));
    LocalMux I__3539 (
            .O(N__24980),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__3538 (
            .O(N__24977),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__3537 (
            .O(N__24974),
            .I(N__24970));
    CascadeMux I__3536 (
            .O(N__24973),
            .I(N__24967));
    InMux I__3535 (
            .O(N__24970),
            .I(N__24964));
    InMux I__3534 (
            .O(N__24967),
            .I(N__24959));
    LocalMux I__3533 (
            .O(N__24964),
            .I(N__24956));
    InMux I__3532 (
            .O(N__24963),
            .I(N__24953));
    InMux I__3531 (
            .O(N__24962),
            .I(N__24950));
    LocalMux I__3530 (
            .O(N__24959),
            .I(N__24943));
    Sp12to4 I__3529 (
            .O(N__24956),
            .I(N__24943));
    LocalMux I__3528 (
            .O(N__24953),
            .I(N__24943));
    LocalMux I__3527 (
            .O(N__24950),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv12 I__3526 (
            .O(N__24943),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__3525 (
            .O(N__24938),
            .I(N__24932));
    InMux I__3524 (
            .O(N__24937),
            .I(N__24932));
    LocalMux I__3523 (
            .O(N__24932),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__3522 (
            .O(N__24929),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    CascadeMux I__3521 (
            .O(N__24926),
            .I(N__24923));
    InMux I__3520 (
            .O(N__24923),
            .I(N__24920));
    LocalMux I__3519 (
            .O(N__24920),
            .I(N__24917));
    Span4Mux_h I__3518 (
            .O(N__24917),
            .I(N__24912));
    InMux I__3517 (
            .O(N__24916),
            .I(N__24908));
    InMux I__3516 (
            .O(N__24915),
            .I(N__24905));
    Span4Mux_v I__3515 (
            .O(N__24912),
            .I(N__24902));
    InMux I__3514 (
            .O(N__24911),
            .I(N__24899));
    LocalMux I__3513 (
            .O(N__24908),
            .I(N__24894));
    LocalMux I__3512 (
            .O(N__24905),
            .I(N__24894));
    Odrv4 I__3511 (
            .O(N__24902),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__3510 (
            .O(N__24899),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__3509 (
            .O(N__24894),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__3508 (
            .O(N__24887),
            .I(N__24881));
    InMux I__3507 (
            .O(N__24886),
            .I(N__24881));
    LocalMux I__3506 (
            .O(N__24881),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__3505 (
            .O(N__24878),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__3504 (
            .O(N__24875),
            .I(N__24872));
    InMux I__3503 (
            .O(N__24872),
            .I(N__24869));
    LocalMux I__3502 (
            .O(N__24869),
            .I(N__24866));
    Span4Mux_h I__3501 (
            .O(N__24866),
            .I(N__24860));
    CascadeMux I__3500 (
            .O(N__24865),
            .I(N__24857));
    InMux I__3499 (
            .O(N__24864),
            .I(N__24854));
    InMux I__3498 (
            .O(N__24863),
            .I(N__24851));
    Span4Mux_v I__3497 (
            .O(N__24860),
            .I(N__24848));
    InMux I__3496 (
            .O(N__24857),
            .I(N__24845));
    LocalMux I__3495 (
            .O(N__24854),
            .I(N__24840));
    LocalMux I__3494 (
            .O(N__24851),
            .I(N__24840));
    Odrv4 I__3493 (
            .O(N__24848),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__3492 (
            .O(N__24845),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__3491 (
            .O(N__24840),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__3490 (
            .O(N__24833),
            .I(N__24827));
    InMux I__3489 (
            .O(N__24832),
            .I(N__24827));
    LocalMux I__3488 (
            .O(N__24827),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__3487 (
            .O(N__24824),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__3486 (
            .O(N__24821),
            .I(N__24818));
    InMux I__3485 (
            .O(N__24818),
            .I(N__24815));
    LocalMux I__3484 (
            .O(N__24815),
            .I(N__24811));
    InMux I__3483 (
            .O(N__24814),
            .I(N__24808));
    Span4Mux_v I__3482 (
            .O(N__24811),
            .I(N__24803));
    LocalMux I__3481 (
            .O(N__24808),
            .I(N__24800));
    InMux I__3480 (
            .O(N__24807),
            .I(N__24795));
    InMux I__3479 (
            .O(N__24806),
            .I(N__24795));
    Odrv4 I__3478 (
            .O(N__24803),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__3477 (
            .O(N__24800),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__3476 (
            .O(N__24795),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__3475 (
            .O(N__24788),
            .I(N__24784));
    InMux I__3474 (
            .O(N__24787),
            .I(N__24779));
    InMux I__3473 (
            .O(N__24784),
            .I(N__24779));
    LocalMux I__3472 (
            .O(N__24779),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__3471 (
            .O(N__24776),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    InMux I__3470 (
            .O(N__24773),
            .I(N__24767));
    InMux I__3469 (
            .O(N__24772),
            .I(N__24767));
    LocalMux I__3468 (
            .O(N__24767),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__3467 (
            .O(N__24764),
            .I(bfn_5_22_0_));
    CascadeMux I__3466 (
            .O(N__24761),
            .I(N__24758));
    InMux I__3465 (
            .O(N__24758),
            .I(N__24754));
    CascadeMux I__3464 (
            .O(N__24757),
            .I(N__24751));
    LocalMux I__3463 (
            .O(N__24754),
            .I(N__24748));
    InMux I__3462 (
            .O(N__24751),
            .I(N__24745));
    Odrv4 I__3461 (
            .O(N__24748),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    LocalMux I__3460 (
            .O(N__24745),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    CascadeMux I__3459 (
            .O(N__24740),
            .I(N__24737));
    InMux I__3458 (
            .O(N__24737),
            .I(N__24734));
    LocalMux I__3457 (
            .O(N__24734),
            .I(N__24730));
    InMux I__3456 (
            .O(N__24733),
            .I(N__24727));
    Span4Mux_h I__3455 (
            .O(N__24730),
            .I(N__24722));
    LocalMux I__3454 (
            .O(N__24727),
            .I(N__24719));
    InMux I__3453 (
            .O(N__24726),
            .I(N__24716));
    InMux I__3452 (
            .O(N__24725),
            .I(N__24713));
    Span4Mux_v I__3451 (
            .O(N__24722),
            .I(N__24710));
    Span4Mux_v I__3450 (
            .O(N__24719),
            .I(N__24707));
    LocalMux I__3449 (
            .O(N__24716),
            .I(N__24704));
    LocalMux I__3448 (
            .O(N__24713),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__3447 (
            .O(N__24710),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__3446 (
            .O(N__24707),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv12 I__3445 (
            .O(N__24704),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__3444 (
            .O(N__24695),
            .I(N__24689));
    InMux I__3443 (
            .O(N__24694),
            .I(N__24689));
    LocalMux I__3442 (
            .O(N__24689),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__3441 (
            .O(N__24686),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    CascadeMux I__3440 (
            .O(N__24683),
            .I(N__24680));
    InMux I__3439 (
            .O(N__24680),
            .I(N__24675));
    InMux I__3438 (
            .O(N__24679),
            .I(N__24672));
    InMux I__3437 (
            .O(N__24678),
            .I(N__24669));
    LocalMux I__3436 (
            .O(N__24675),
            .I(N__24663));
    LocalMux I__3435 (
            .O(N__24672),
            .I(N__24663));
    LocalMux I__3434 (
            .O(N__24669),
            .I(N__24660));
    CascadeMux I__3433 (
            .O(N__24668),
            .I(N__24657));
    Span4Mux_v I__3432 (
            .O(N__24663),
            .I(N__24654));
    Span4Mux_v I__3431 (
            .O(N__24660),
            .I(N__24651));
    InMux I__3430 (
            .O(N__24657),
            .I(N__24648));
    Odrv4 I__3429 (
            .O(N__24654),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__3428 (
            .O(N__24651),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__3427 (
            .O(N__24648),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__3426 (
            .O(N__24641),
            .I(N__24635));
    InMux I__3425 (
            .O(N__24640),
            .I(N__24635));
    LocalMux I__3424 (
            .O(N__24635),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__3423 (
            .O(N__24632),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    CascadeMux I__3422 (
            .O(N__24629),
            .I(N__24624));
    InMux I__3421 (
            .O(N__24628),
            .I(N__24621));
    InMux I__3420 (
            .O(N__24627),
            .I(N__24618));
    InMux I__3419 (
            .O(N__24624),
            .I(N__24615));
    LocalMux I__3418 (
            .O(N__24621),
            .I(N__24609));
    LocalMux I__3417 (
            .O(N__24618),
            .I(N__24609));
    LocalMux I__3416 (
            .O(N__24615),
            .I(N__24606));
    InMux I__3415 (
            .O(N__24614),
            .I(N__24603));
    Span4Mux_v I__3414 (
            .O(N__24609),
            .I(N__24600));
    Odrv12 I__3413 (
            .O(N__24606),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__3412 (
            .O(N__24603),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__3411 (
            .O(N__24600),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__3410 (
            .O(N__24593),
            .I(N__24589));
    InMux I__3409 (
            .O(N__24592),
            .I(N__24586));
    InMux I__3408 (
            .O(N__24589),
            .I(N__24583));
    LocalMux I__3407 (
            .O(N__24586),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    LocalMux I__3406 (
            .O(N__24583),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__3405 (
            .O(N__24578),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__3404 (
            .O(N__24575),
            .I(N__24572));
    InMux I__3403 (
            .O(N__24572),
            .I(N__24568));
    CascadeMux I__3402 (
            .O(N__24571),
            .I(N__24565));
    LocalMux I__3401 (
            .O(N__24568),
            .I(N__24561));
    InMux I__3400 (
            .O(N__24565),
            .I(N__24558));
    InMux I__3399 (
            .O(N__24564),
            .I(N__24555));
    Span4Mux_v I__3398 (
            .O(N__24561),
            .I(N__24552));
    LocalMux I__3397 (
            .O(N__24558),
            .I(N__24548));
    LocalMux I__3396 (
            .O(N__24555),
            .I(N__24545));
    Span4Mux_v I__3395 (
            .O(N__24552),
            .I(N__24542));
    InMux I__3394 (
            .O(N__24551),
            .I(N__24539));
    Span4Mux_s3_h I__3393 (
            .O(N__24548),
            .I(N__24534));
    Span4Mux_v I__3392 (
            .O(N__24545),
            .I(N__24534));
    Odrv4 I__3391 (
            .O(N__24542),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__3390 (
            .O(N__24539),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__3389 (
            .O(N__24534),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__3388 (
            .O(N__24527),
            .I(N__24521));
    InMux I__3387 (
            .O(N__24526),
            .I(N__24521));
    LocalMux I__3386 (
            .O(N__24521),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__3385 (
            .O(N__24518),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    CascadeMux I__3384 (
            .O(N__24515),
            .I(N__24512));
    InMux I__3383 (
            .O(N__24512),
            .I(N__24509));
    LocalMux I__3382 (
            .O(N__24509),
            .I(N__24505));
    CascadeMux I__3381 (
            .O(N__24508),
            .I(N__24502));
    Span4Mux_h I__3380 (
            .O(N__24505),
            .I(N__24497));
    InMux I__3379 (
            .O(N__24502),
            .I(N__24494));
    InMux I__3378 (
            .O(N__24501),
            .I(N__24491));
    CascadeMux I__3377 (
            .O(N__24500),
            .I(N__24488));
    Span4Mux_h I__3376 (
            .O(N__24497),
            .I(N__24481));
    LocalMux I__3375 (
            .O(N__24494),
            .I(N__24481));
    LocalMux I__3374 (
            .O(N__24491),
            .I(N__24481));
    InMux I__3373 (
            .O(N__24488),
            .I(N__24478));
    Span4Mux_v I__3372 (
            .O(N__24481),
            .I(N__24475));
    LocalMux I__3371 (
            .O(N__24478),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__3370 (
            .O(N__24475),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__3369 (
            .O(N__24470),
            .I(N__24464));
    InMux I__3368 (
            .O(N__24469),
            .I(N__24464));
    LocalMux I__3367 (
            .O(N__24464),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__3366 (
            .O(N__24461),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__3365 (
            .O(N__24458),
            .I(N__24455));
    LocalMux I__3364 (
            .O(N__24455),
            .I(N__24450));
    InMux I__3363 (
            .O(N__24454),
            .I(N__24447));
    InMux I__3362 (
            .O(N__24453),
            .I(N__24443));
    Span4Mux_v I__3361 (
            .O(N__24450),
            .I(N__24438));
    LocalMux I__3360 (
            .O(N__24447),
            .I(N__24438));
    InMux I__3359 (
            .O(N__24446),
            .I(N__24435));
    LocalMux I__3358 (
            .O(N__24443),
            .I(N__24430));
    Span4Mux_h I__3357 (
            .O(N__24438),
            .I(N__24430));
    LocalMux I__3356 (
            .O(N__24435),
            .I(N__24427));
    Span4Mux_v I__3355 (
            .O(N__24430),
            .I(N__24424));
    Odrv12 I__3354 (
            .O(N__24427),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__3353 (
            .O(N__24424),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__3352 (
            .O(N__24419),
            .I(N__24415));
    InMux I__3351 (
            .O(N__24418),
            .I(N__24410));
    InMux I__3350 (
            .O(N__24415),
            .I(N__24410));
    LocalMux I__3349 (
            .O(N__24410),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__3348 (
            .O(N__24407),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    CascadeMux I__3347 (
            .O(N__24404),
            .I(N__24401));
    InMux I__3346 (
            .O(N__24401),
            .I(N__24397));
    CascadeMux I__3345 (
            .O(N__24400),
            .I(N__24393));
    LocalMux I__3344 (
            .O(N__24397),
            .I(N__24389));
    InMux I__3343 (
            .O(N__24396),
            .I(N__24386));
    InMux I__3342 (
            .O(N__24393),
            .I(N__24383));
    InMux I__3341 (
            .O(N__24392),
            .I(N__24380));
    Span4Mux_v I__3340 (
            .O(N__24389),
            .I(N__24377));
    LocalMux I__3339 (
            .O(N__24386),
            .I(N__24374));
    LocalMux I__3338 (
            .O(N__24383),
            .I(N__24369));
    LocalMux I__3337 (
            .O(N__24380),
            .I(N__24369));
    Odrv4 I__3336 (
            .O(N__24377),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__3335 (
            .O(N__24374),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__3334 (
            .O(N__24369),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    CascadeMux I__3333 (
            .O(N__24362),
            .I(N__24359));
    InMux I__3332 (
            .O(N__24359),
            .I(N__24355));
    InMux I__3331 (
            .O(N__24358),
            .I(N__24352));
    LocalMux I__3330 (
            .O(N__24355),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    LocalMux I__3329 (
            .O(N__24352),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__3328 (
            .O(N__24347),
            .I(bfn_5_21_0_));
    CascadeMux I__3327 (
            .O(N__24344),
            .I(N__24341));
    InMux I__3326 (
            .O(N__24341),
            .I(N__24338));
    LocalMux I__3325 (
            .O(N__24338),
            .I(N__24334));
    InMux I__3324 (
            .O(N__24337),
            .I(N__24330));
    Span4Mux_h I__3323 (
            .O(N__24334),
            .I(N__24326));
    InMux I__3322 (
            .O(N__24333),
            .I(N__24323));
    LocalMux I__3321 (
            .O(N__24330),
            .I(N__24320));
    InMux I__3320 (
            .O(N__24329),
            .I(N__24317));
    Span4Mux_v I__3319 (
            .O(N__24326),
            .I(N__24310));
    LocalMux I__3318 (
            .O(N__24323),
            .I(N__24310));
    Span4Mux_v I__3317 (
            .O(N__24320),
            .I(N__24310));
    LocalMux I__3316 (
            .O(N__24317),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__3315 (
            .O(N__24310),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__3314 (
            .O(N__24305),
            .I(N__24301));
    InMux I__3313 (
            .O(N__24304),
            .I(N__24298));
    LocalMux I__3312 (
            .O(N__24301),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__3311 (
            .O(N__24298),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__3310 (
            .O(N__24293),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__3309 (
            .O(N__24290),
            .I(N__24287));
    LocalMux I__3308 (
            .O(N__24287),
            .I(N__24284));
    Odrv12 I__3307 (
            .O(N__24284),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__3306 (
            .O(N__24281),
            .I(N__24278));
    InMux I__3305 (
            .O(N__24278),
            .I(N__24273));
    InMux I__3304 (
            .O(N__24277),
            .I(N__24270));
    InMux I__3303 (
            .O(N__24276),
            .I(N__24267));
    LocalMux I__3302 (
            .O(N__24273),
            .I(N__24264));
    LocalMux I__3301 (
            .O(N__24270),
            .I(N__24261));
    LocalMux I__3300 (
            .O(N__24267),
            .I(N__24256));
    Span4Mux_h I__3299 (
            .O(N__24264),
            .I(N__24256));
    Span4Mux_v I__3298 (
            .O(N__24261),
            .I(N__24252));
    Span4Mux_v I__3297 (
            .O(N__24256),
            .I(N__24249));
    InMux I__3296 (
            .O(N__24255),
            .I(N__24246));
    Odrv4 I__3295 (
            .O(N__24252),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3294 (
            .O(N__24249),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__3293 (
            .O(N__24246),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__3292 (
            .O(N__24239),
            .I(N__24234));
    InMux I__3291 (
            .O(N__24238),
            .I(N__24229));
    InMux I__3290 (
            .O(N__24237),
            .I(N__24229));
    LocalMux I__3289 (
            .O(N__24234),
            .I(N__24224));
    LocalMux I__3288 (
            .O(N__24229),
            .I(N__24224));
    Span4Mux_v I__3287 (
            .O(N__24224),
            .I(N__24221));
    Odrv4 I__3286 (
            .O(N__24221),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__3285 (
            .O(N__24218),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__3284 (
            .O(N__24215),
            .I(N__24212));
    LocalMux I__3283 (
            .O(N__24212),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__3282 (
            .O(N__24209),
            .I(N__24204));
    CascadeMux I__3281 (
            .O(N__24208),
            .I(N__24201));
    CascadeMux I__3280 (
            .O(N__24207),
            .I(N__24198));
    InMux I__3279 (
            .O(N__24204),
            .I(N__24194));
    InMux I__3278 (
            .O(N__24201),
            .I(N__24191));
    InMux I__3277 (
            .O(N__24198),
            .I(N__24188));
    InMux I__3276 (
            .O(N__24197),
            .I(N__24185));
    LocalMux I__3275 (
            .O(N__24194),
            .I(N__24182));
    LocalMux I__3274 (
            .O(N__24191),
            .I(N__24179));
    LocalMux I__3273 (
            .O(N__24188),
            .I(N__24176));
    LocalMux I__3272 (
            .O(N__24185),
            .I(N__24173));
    Span4Mux_v I__3271 (
            .O(N__24182),
            .I(N__24170));
    Span4Mux_h I__3270 (
            .O(N__24179),
            .I(N__24167));
    Odrv4 I__3269 (
            .O(N__24176),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__3268 (
            .O(N__24173),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__3267 (
            .O(N__24170),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__3266 (
            .O(N__24167),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__3265 (
            .O(N__24158),
            .I(N__24152));
    InMux I__3264 (
            .O(N__24157),
            .I(N__24149));
    InMux I__3263 (
            .O(N__24156),
            .I(N__24144));
    InMux I__3262 (
            .O(N__24155),
            .I(N__24144));
    LocalMux I__3261 (
            .O(N__24152),
            .I(N__24139));
    LocalMux I__3260 (
            .O(N__24149),
            .I(N__24139));
    LocalMux I__3259 (
            .O(N__24144),
            .I(N__24136));
    Span4Mux_v I__3258 (
            .O(N__24139),
            .I(N__24133));
    Span4Mux_h I__3257 (
            .O(N__24136),
            .I(N__24130));
    Odrv4 I__3256 (
            .O(N__24133),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__3255 (
            .O(N__24130),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__3254 (
            .O(N__24125),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__3253 (
            .O(N__24122),
            .I(N__24119));
    LocalMux I__3252 (
            .O(N__24119),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__3251 (
            .O(N__24116),
            .I(N__24112));
    InMux I__3250 (
            .O(N__24115),
            .I(N__24108));
    InMux I__3249 (
            .O(N__24112),
            .I(N__24105));
    InMux I__3248 (
            .O(N__24111),
            .I(N__24101));
    LocalMux I__3247 (
            .O(N__24108),
            .I(N__24098));
    LocalMux I__3246 (
            .O(N__24105),
            .I(N__24095));
    InMux I__3245 (
            .O(N__24104),
            .I(N__24092));
    LocalMux I__3244 (
            .O(N__24101),
            .I(N__24089));
    Span4Mux_v I__3243 (
            .O(N__24098),
            .I(N__24086));
    Span12Mux_h I__3242 (
            .O(N__24095),
            .I(N__24081));
    LocalMux I__3241 (
            .O(N__24092),
            .I(N__24081));
    Span4Mux_h I__3240 (
            .O(N__24089),
            .I(N__24078));
    Odrv4 I__3239 (
            .O(N__24086),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv12 I__3238 (
            .O(N__24081),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__3237 (
            .O(N__24078),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    CascadeMux I__3236 (
            .O(N__24071),
            .I(N__24067));
    InMux I__3235 (
            .O(N__24070),
            .I(N__24063));
    InMux I__3234 (
            .O(N__24067),
            .I(N__24060));
    InMux I__3233 (
            .O(N__24066),
            .I(N__24057));
    LocalMux I__3232 (
            .O(N__24063),
            .I(N__24054));
    LocalMux I__3231 (
            .O(N__24060),
            .I(N__24051));
    LocalMux I__3230 (
            .O(N__24057),
            .I(N__24048));
    Span4Mux_v I__3229 (
            .O(N__24054),
            .I(N__24045));
    Span4Mux_h I__3228 (
            .O(N__24051),
            .I(N__24042));
    Span4Mux_h I__3227 (
            .O(N__24048),
            .I(N__24039));
    Odrv4 I__3226 (
            .O(N__24045),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__3225 (
            .O(N__24042),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__3224 (
            .O(N__24039),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__3223 (
            .O(N__24032),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__3222 (
            .O(N__24029),
            .I(N__24025));
    CascadeMux I__3221 (
            .O(N__24028),
            .I(N__24021));
    LocalMux I__3220 (
            .O(N__24025),
            .I(N__24018));
    InMux I__3219 (
            .O(N__24024),
            .I(N__24015));
    InMux I__3218 (
            .O(N__24021),
            .I(N__24012));
    Span4Mux_v I__3217 (
            .O(N__24018),
            .I(N__24007));
    LocalMux I__3216 (
            .O(N__24015),
            .I(N__24007));
    LocalMux I__3215 (
            .O(N__24012),
            .I(N__24004));
    Span4Mux_v I__3214 (
            .O(N__24007),
            .I(N__23998));
    Span4Mux_h I__3213 (
            .O(N__24004),
            .I(N__23998));
    InMux I__3212 (
            .O(N__24003),
            .I(N__23995));
    Span4Mux_v I__3211 (
            .O(N__23998),
            .I(N__23992));
    LocalMux I__3210 (
            .O(N__23995),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__3209 (
            .O(N__23992),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__3208 (
            .O(N__23987),
            .I(N__23984));
    InMux I__3207 (
            .O(N__23984),
            .I(N__23981));
    LocalMux I__3206 (
            .O(N__23981),
            .I(N__23978));
    Odrv4 I__3205 (
            .O(N__23978),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__3204 (
            .O(N__23975),
            .I(N__23970));
    InMux I__3203 (
            .O(N__23974),
            .I(N__23965));
    InMux I__3202 (
            .O(N__23973),
            .I(N__23965));
    LocalMux I__3201 (
            .O(N__23970),
            .I(N__23962));
    LocalMux I__3200 (
            .O(N__23965),
            .I(N__23959));
    Span4Mux_v I__3199 (
            .O(N__23962),
            .I(N__23956));
    Span4Mux_h I__3198 (
            .O(N__23959),
            .I(N__23953));
    Odrv4 I__3197 (
            .O(N__23956),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__3196 (
            .O(N__23953),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__3195 (
            .O(N__23948),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__3194 (
            .O(N__23945),
            .I(N__23942));
    LocalMux I__3193 (
            .O(N__23942),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__3192 (
            .O(N__23939),
            .I(N__23936));
    InMux I__3191 (
            .O(N__23936),
            .I(N__23933));
    LocalMux I__3190 (
            .O(N__23933),
            .I(N__23928));
    InMux I__3189 (
            .O(N__23932),
            .I(N__23925));
    InMux I__3188 (
            .O(N__23931),
            .I(N__23922));
    Span4Mux_h I__3187 (
            .O(N__23928),
            .I(N__23914));
    LocalMux I__3186 (
            .O(N__23925),
            .I(N__23914));
    LocalMux I__3185 (
            .O(N__23922),
            .I(N__23914));
    InMux I__3184 (
            .O(N__23921),
            .I(N__23911));
    Span4Mux_v I__3183 (
            .O(N__23914),
            .I(N__23908));
    LocalMux I__3182 (
            .O(N__23911),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__3181 (
            .O(N__23908),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__3180 (
            .O(N__23903),
            .I(N__23898));
    InMux I__3179 (
            .O(N__23902),
            .I(N__23895));
    InMux I__3178 (
            .O(N__23901),
            .I(N__23892));
    LocalMux I__3177 (
            .O(N__23898),
            .I(N__23889));
    LocalMux I__3176 (
            .O(N__23895),
            .I(N__23886));
    LocalMux I__3175 (
            .O(N__23892),
            .I(N__23883));
    Span4Mux_v I__3174 (
            .O(N__23889),
            .I(N__23880));
    Span4Mux_h I__3173 (
            .O(N__23886),
            .I(N__23877));
    Span4Mux_h I__3172 (
            .O(N__23883),
            .I(N__23874));
    Odrv4 I__3171 (
            .O(N__23880),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__3170 (
            .O(N__23877),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__3169 (
            .O(N__23874),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__3168 (
            .O(N__23867),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__3167 (
            .O(N__23864),
            .I(N__23861));
    LocalMux I__3166 (
            .O(N__23861),
            .I(N__23858));
    Odrv4 I__3165 (
            .O(N__23858),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__3164 (
            .O(N__23855),
            .I(N__23852));
    InMux I__3163 (
            .O(N__23852),
            .I(N__23849));
    LocalMux I__3162 (
            .O(N__23849),
            .I(N__23844));
    InMux I__3161 (
            .O(N__23848),
            .I(N__23841));
    InMux I__3160 (
            .O(N__23847),
            .I(N__23838));
    Span4Mux_v I__3159 (
            .O(N__23844),
            .I(N__23835));
    LocalMux I__3158 (
            .O(N__23841),
            .I(N__23829));
    LocalMux I__3157 (
            .O(N__23838),
            .I(N__23829));
    Span4Mux_v I__3156 (
            .O(N__23835),
            .I(N__23826));
    InMux I__3155 (
            .O(N__23834),
            .I(N__23823));
    Span4Mux_v I__3154 (
            .O(N__23829),
            .I(N__23820));
    Odrv4 I__3153 (
            .O(N__23826),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3152 (
            .O(N__23823),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__3151 (
            .O(N__23820),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__3150 (
            .O(N__23813),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    CascadeMux I__3149 (
            .O(N__23810),
            .I(N__23807));
    InMux I__3148 (
            .O(N__23807),
            .I(N__23803));
    InMux I__3147 (
            .O(N__23806),
            .I(N__23800));
    LocalMux I__3146 (
            .O(N__23803),
            .I(N__23797));
    LocalMux I__3145 (
            .O(N__23800),
            .I(N__23793));
    Span4Mux_h I__3144 (
            .O(N__23797),
            .I(N__23790));
    InMux I__3143 (
            .O(N__23796),
            .I(N__23786));
    Span4Mux_v I__3142 (
            .O(N__23793),
            .I(N__23783));
    Span4Mux_v I__3141 (
            .O(N__23790),
            .I(N__23780));
    InMux I__3140 (
            .O(N__23789),
            .I(N__23777));
    LocalMux I__3139 (
            .O(N__23786),
            .I(N__23774));
    Odrv4 I__3138 (
            .O(N__23783),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__3137 (
            .O(N__23780),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__3136 (
            .O(N__23777),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__3135 (
            .O(N__23774),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__3134 (
            .O(N__23765),
            .I(bfn_5_20_0_));
    CascadeMux I__3133 (
            .O(N__23762),
            .I(N__23758));
    CascadeMux I__3132 (
            .O(N__23761),
            .I(N__23754));
    InMux I__3131 (
            .O(N__23758),
            .I(N__23751));
    InMux I__3130 (
            .O(N__23757),
            .I(N__23748));
    InMux I__3129 (
            .O(N__23754),
            .I(N__23745));
    LocalMux I__3128 (
            .O(N__23751),
            .I(N__23742));
    LocalMux I__3127 (
            .O(N__23748),
            .I(N__23737));
    LocalMux I__3126 (
            .O(N__23745),
            .I(N__23737));
    Span4Mux_v I__3125 (
            .O(N__23742),
            .I(N__23731));
    Span4Mux_v I__3124 (
            .O(N__23737),
            .I(N__23731));
    InMux I__3123 (
            .O(N__23736),
            .I(N__23728));
    Odrv4 I__3122 (
            .O(N__23731),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__3121 (
            .O(N__23728),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__3120 (
            .O(N__23723),
            .I(N__23717));
    InMux I__3119 (
            .O(N__23722),
            .I(N__23717));
    LocalMux I__3118 (
            .O(N__23717),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__3117 (
            .O(N__23714),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    CascadeMux I__3116 (
            .O(N__23711),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ));
    InMux I__3115 (
            .O(N__23708),
            .I(N__23705));
    LocalMux I__3114 (
            .O(N__23705),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__3113 (
            .O(N__23702),
            .I(N__23699));
    LocalMux I__3112 (
            .O(N__23699),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ));
    InMux I__3111 (
            .O(N__23696),
            .I(N__23693));
    LocalMux I__3110 (
            .O(N__23693),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__3109 (
            .O(N__23690),
            .I(N__23686));
    InMux I__3108 (
            .O(N__23689),
            .I(N__23683));
    LocalMux I__3107 (
            .O(N__23686),
            .I(N__23678));
    LocalMux I__3106 (
            .O(N__23683),
            .I(N__23678));
    Odrv4 I__3105 (
            .O(N__23678),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__3104 (
            .O(N__23675),
            .I(N__23670));
    InMux I__3103 (
            .O(N__23674),
            .I(N__23667));
    InMux I__3102 (
            .O(N__23673),
            .I(N__23664));
    InMux I__3101 (
            .O(N__23670),
            .I(N__23661));
    LocalMux I__3100 (
            .O(N__23667),
            .I(N__23655));
    LocalMux I__3099 (
            .O(N__23664),
            .I(N__23655));
    LocalMux I__3098 (
            .O(N__23661),
            .I(N__23652));
    InMux I__3097 (
            .O(N__23660),
            .I(N__23648));
    Span4Mux_v I__3096 (
            .O(N__23655),
            .I(N__23645));
    Span12Mux_h I__3095 (
            .O(N__23652),
            .I(N__23642));
    InMux I__3094 (
            .O(N__23651),
            .I(N__23639));
    LocalMux I__3093 (
            .O(N__23648),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__3092 (
            .O(N__23645),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__3091 (
            .O(N__23642),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__3090 (
            .O(N__23639),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__3089 (
            .O(N__23630),
            .I(N__23627));
    LocalMux I__3088 (
            .O(N__23627),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__3087 (
            .O(N__23624),
            .I(N__23620));
    InMux I__3086 (
            .O(N__23623),
            .I(N__23617));
    InMux I__3085 (
            .O(N__23620),
            .I(N__23614));
    LocalMux I__3084 (
            .O(N__23617),
            .I(N__23608));
    LocalMux I__3083 (
            .O(N__23614),
            .I(N__23608));
    CascadeMux I__3082 (
            .O(N__23613),
            .I(N__23605));
    Sp12to4 I__3081 (
            .O(N__23608),
            .I(N__23602));
    InMux I__3080 (
            .O(N__23605),
            .I(N__23599));
    Odrv12 I__3079 (
            .O(N__23602),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__3078 (
            .O(N__23599),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__3077 (
            .O(N__23594),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__3076 (
            .O(N__23591),
            .I(N__23588));
    LocalMux I__3075 (
            .O(N__23588),
            .I(N__23585));
    Span12Mux_v I__3074 (
            .O(N__23585),
            .I(N__23582));
    Span12Mux_h I__3073 (
            .O(N__23582),
            .I(N__23579));
    Odrv12 I__3072 (
            .O(N__23579),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    CascadeMux I__3071 (
            .O(N__23576),
            .I(N__23573));
    InMux I__3070 (
            .O(N__23573),
            .I(N__23570));
    LocalMux I__3069 (
            .O(N__23570),
            .I(N__23567));
    Odrv4 I__3068 (
            .O(N__23567),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__3067 (
            .O(N__23564),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__3066 (
            .O(N__23561),
            .I(N__23558));
    LocalMux I__3065 (
            .O(N__23558),
            .I(N__23555));
    Span4Mux_v I__3064 (
            .O(N__23555),
            .I(N__23552));
    Sp12to4 I__3063 (
            .O(N__23552),
            .I(N__23549));
    Span12Mux_h I__3062 (
            .O(N__23549),
            .I(N__23546));
    Span12Mux_h I__3061 (
            .O(N__23546),
            .I(N__23543));
    Odrv12 I__3060 (
            .O(N__23543),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    CascadeMux I__3059 (
            .O(N__23540),
            .I(N__23537));
    InMux I__3058 (
            .O(N__23537),
            .I(N__23534));
    LocalMux I__3057 (
            .O(N__23534),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__3056 (
            .O(N__23531),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__3055 (
            .O(N__23528),
            .I(N__23525));
    LocalMux I__3054 (
            .O(N__23525),
            .I(N__23522));
    Span4Mux_v I__3053 (
            .O(N__23522),
            .I(N__23519));
    Sp12to4 I__3052 (
            .O(N__23519),
            .I(N__23516));
    Span12Mux_h I__3051 (
            .O(N__23516),
            .I(N__23513));
    Span12Mux_h I__3050 (
            .O(N__23513),
            .I(N__23510));
    Odrv12 I__3049 (
            .O(N__23510),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    CascadeMux I__3048 (
            .O(N__23507),
            .I(N__23504));
    InMux I__3047 (
            .O(N__23504),
            .I(N__23501));
    LocalMux I__3046 (
            .O(N__23501),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__3045 (
            .O(N__23498),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__3044 (
            .O(N__23495),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    CascadeMux I__3043 (
            .O(N__23492),
            .I(N__23489));
    InMux I__3042 (
            .O(N__23489),
            .I(N__23486));
    LocalMux I__3041 (
            .O(N__23486),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    InMux I__3040 (
            .O(N__23483),
            .I(N__23480));
    LocalMux I__3039 (
            .O(N__23480),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    CascadeMux I__3038 (
            .O(N__23477),
            .I(N__23463));
    CascadeMux I__3037 (
            .O(N__23476),
            .I(N__23460));
    CascadeMux I__3036 (
            .O(N__23475),
            .I(N__23457));
    CascadeMux I__3035 (
            .O(N__23474),
            .I(N__23454));
    CascadeMux I__3034 (
            .O(N__23473),
            .I(N__23450));
    CascadeMux I__3033 (
            .O(N__23472),
            .I(N__23447));
    CascadeMux I__3032 (
            .O(N__23471),
            .I(N__23444));
    CascadeMux I__3031 (
            .O(N__23470),
            .I(N__23441));
    InMux I__3030 (
            .O(N__23469),
            .I(N__23431));
    InMux I__3029 (
            .O(N__23468),
            .I(N__23431));
    InMux I__3028 (
            .O(N__23467),
            .I(N__23417));
    InMux I__3027 (
            .O(N__23466),
            .I(N__23410));
    InMux I__3026 (
            .O(N__23463),
            .I(N__23410));
    InMux I__3025 (
            .O(N__23460),
            .I(N__23410));
    InMux I__3024 (
            .O(N__23457),
            .I(N__23403));
    InMux I__3023 (
            .O(N__23454),
            .I(N__23403));
    InMux I__3022 (
            .O(N__23453),
            .I(N__23403));
    InMux I__3021 (
            .O(N__23450),
            .I(N__23390));
    InMux I__3020 (
            .O(N__23447),
            .I(N__23390));
    InMux I__3019 (
            .O(N__23444),
            .I(N__23390));
    InMux I__3018 (
            .O(N__23441),
            .I(N__23390));
    InMux I__3017 (
            .O(N__23440),
            .I(N__23390));
    InMux I__3016 (
            .O(N__23439),
            .I(N__23390));
    InMux I__3015 (
            .O(N__23438),
            .I(N__23387));
    InMux I__3014 (
            .O(N__23437),
            .I(N__23380));
    InMux I__3013 (
            .O(N__23436),
            .I(N__23380));
    LocalMux I__3012 (
            .O(N__23431),
            .I(N__23377));
    InMux I__3011 (
            .O(N__23430),
            .I(N__23362));
    InMux I__3010 (
            .O(N__23429),
            .I(N__23362));
    InMux I__3009 (
            .O(N__23428),
            .I(N__23362));
    InMux I__3008 (
            .O(N__23427),
            .I(N__23362));
    InMux I__3007 (
            .O(N__23426),
            .I(N__23362));
    InMux I__3006 (
            .O(N__23425),
            .I(N__23362));
    InMux I__3005 (
            .O(N__23424),
            .I(N__23362));
    InMux I__3004 (
            .O(N__23423),
            .I(N__23353));
    InMux I__3003 (
            .O(N__23422),
            .I(N__23353));
    InMux I__3002 (
            .O(N__23421),
            .I(N__23353));
    InMux I__3001 (
            .O(N__23420),
            .I(N__23353));
    LocalMux I__3000 (
            .O(N__23417),
            .I(N__23350));
    LocalMux I__2999 (
            .O(N__23410),
            .I(N__23345));
    LocalMux I__2998 (
            .O(N__23403),
            .I(N__23345));
    LocalMux I__2997 (
            .O(N__23390),
            .I(N__23340));
    LocalMux I__2996 (
            .O(N__23387),
            .I(N__23340));
    InMux I__2995 (
            .O(N__23386),
            .I(N__23335));
    InMux I__2994 (
            .O(N__23385),
            .I(N__23335));
    LocalMux I__2993 (
            .O(N__23380),
            .I(N__23330));
    Span4Mux_h I__2992 (
            .O(N__23377),
            .I(N__23330));
    LocalMux I__2991 (
            .O(N__23362),
            .I(N__23321));
    LocalMux I__2990 (
            .O(N__23353),
            .I(N__23321));
    Span4Mux_h I__2989 (
            .O(N__23350),
            .I(N__23321));
    Span4Mux_v I__2988 (
            .O(N__23345),
            .I(N__23321));
    Span4Mux_v I__2987 (
            .O(N__23340),
            .I(N__23318));
    LocalMux I__2986 (
            .O(N__23335),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2985 (
            .O(N__23330),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2984 (
            .O(N__23321),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2983 (
            .O(N__23318),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    InMux I__2982 (
            .O(N__23309),
            .I(N__23306));
    LocalMux I__2981 (
            .O(N__23306),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__2980 (
            .O(N__23303),
            .I(N__23300));
    LocalMux I__2979 (
            .O(N__23300),
            .I(N__23297));
    Span4Mux_h I__2978 (
            .O(N__23297),
            .I(N__23294));
    Odrv4 I__2977 (
            .O(N__23294),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    InMux I__2976 (
            .O(N__23291),
            .I(N__23288));
    LocalMux I__2975 (
            .O(N__23288),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    CascadeMux I__2974 (
            .O(N__23285),
            .I(N__23265));
    CascadeMux I__2973 (
            .O(N__23284),
            .I(N__23259));
    InMux I__2972 (
            .O(N__23283),
            .I(N__23245));
    InMux I__2971 (
            .O(N__23282),
            .I(N__23245));
    InMux I__2970 (
            .O(N__23281),
            .I(N__23245));
    InMux I__2969 (
            .O(N__23280),
            .I(N__23245));
    InMux I__2968 (
            .O(N__23279),
            .I(N__23245));
    InMux I__2967 (
            .O(N__23278),
            .I(N__23245));
    InMux I__2966 (
            .O(N__23277),
            .I(N__23240));
    InMux I__2965 (
            .O(N__23276),
            .I(N__23240));
    InMux I__2964 (
            .O(N__23275),
            .I(N__23233));
    InMux I__2963 (
            .O(N__23274),
            .I(N__23233));
    InMux I__2962 (
            .O(N__23273),
            .I(N__23233));
    InMux I__2961 (
            .O(N__23272),
            .I(N__23226));
    InMux I__2960 (
            .O(N__23271),
            .I(N__23226));
    InMux I__2959 (
            .O(N__23270),
            .I(N__23226));
    InMux I__2958 (
            .O(N__23269),
            .I(N__23217));
    InMux I__2957 (
            .O(N__23268),
            .I(N__23214));
    InMux I__2956 (
            .O(N__23265),
            .I(N__23209));
    InMux I__2955 (
            .O(N__23264),
            .I(N__23209));
    InMux I__2954 (
            .O(N__23263),
            .I(N__23200));
    InMux I__2953 (
            .O(N__23262),
            .I(N__23200));
    InMux I__2952 (
            .O(N__23259),
            .I(N__23200));
    InMux I__2951 (
            .O(N__23258),
            .I(N__23200));
    LocalMux I__2950 (
            .O(N__23245),
            .I(N__23197));
    LocalMux I__2949 (
            .O(N__23240),
            .I(N__23192));
    LocalMux I__2948 (
            .O(N__23233),
            .I(N__23192));
    LocalMux I__2947 (
            .O(N__23226),
            .I(N__23189));
    CascadeMux I__2946 (
            .O(N__23225),
            .I(N__23186));
    CascadeMux I__2945 (
            .O(N__23224),
            .I(N__23183));
    CascadeMux I__2944 (
            .O(N__23223),
            .I(N__23178));
    CascadeMux I__2943 (
            .O(N__23222),
            .I(N__23175));
    CascadeMux I__2942 (
            .O(N__23221),
            .I(N__23172));
    CascadeMux I__2941 (
            .O(N__23220),
            .I(N__23169));
    LocalMux I__2940 (
            .O(N__23217),
            .I(N__23165));
    LocalMux I__2939 (
            .O(N__23214),
            .I(N__23162));
    LocalMux I__2938 (
            .O(N__23209),
            .I(N__23159));
    LocalMux I__2937 (
            .O(N__23200),
            .I(N__23150));
    Span4Mux_h I__2936 (
            .O(N__23197),
            .I(N__23150));
    Span4Mux_h I__2935 (
            .O(N__23192),
            .I(N__23150));
    Span4Mux_v I__2934 (
            .O(N__23189),
            .I(N__23150));
    InMux I__2933 (
            .O(N__23186),
            .I(N__23145));
    InMux I__2932 (
            .O(N__23183),
            .I(N__23145));
    InMux I__2931 (
            .O(N__23182),
            .I(N__23130));
    InMux I__2930 (
            .O(N__23181),
            .I(N__23130));
    InMux I__2929 (
            .O(N__23178),
            .I(N__23130));
    InMux I__2928 (
            .O(N__23175),
            .I(N__23130));
    InMux I__2927 (
            .O(N__23172),
            .I(N__23130));
    InMux I__2926 (
            .O(N__23169),
            .I(N__23130));
    InMux I__2925 (
            .O(N__23168),
            .I(N__23130));
    Span4Mux_h I__2924 (
            .O(N__23165),
            .I(N__23127));
    Span4Mux_v I__2923 (
            .O(N__23162),
            .I(N__23124));
    Span4Mux_v I__2922 (
            .O(N__23159),
            .I(N__23119));
    Span4Mux_v I__2921 (
            .O(N__23150),
            .I(N__23119));
    LocalMux I__2920 (
            .O(N__23145),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__2919 (
            .O(N__23130),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2918 (
            .O(N__23127),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2917 (
            .O(N__23124),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2916 (
            .O(N__23119),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    InMux I__2915 (
            .O(N__23108),
            .I(N__23105));
    LocalMux I__2914 (
            .O(N__23105),
            .I(N__23102));
    Span12Mux_v I__2913 (
            .O(N__23102),
            .I(N__23099));
    Span12Mux_h I__2912 (
            .O(N__23099),
            .I(N__23096));
    Odrv12 I__2911 (
            .O(N__23096),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    CascadeMux I__2910 (
            .O(N__23093),
            .I(N__23090));
    InMux I__2909 (
            .O(N__23090),
            .I(N__23087));
    LocalMux I__2908 (
            .O(N__23087),
            .I(N__23084));
    Odrv4 I__2907 (
            .O(N__23084),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__2906 (
            .O(N__23081),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    InMux I__2905 (
            .O(N__23078),
            .I(N__23075));
    LocalMux I__2904 (
            .O(N__23075),
            .I(N__23072));
    Span4Mux_h I__2903 (
            .O(N__23072),
            .I(N__23069));
    Sp12to4 I__2902 (
            .O(N__23069),
            .I(N__23066));
    Span12Mux_v I__2901 (
            .O(N__23066),
            .I(N__23063));
    Span12Mux_h I__2900 (
            .O(N__23063),
            .I(N__23060));
    Odrv12 I__2899 (
            .O(N__23060),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    CascadeMux I__2898 (
            .O(N__23057),
            .I(N__23054));
    InMux I__2897 (
            .O(N__23054),
            .I(N__23051));
    LocalMux I__2896 (
            .O(N__23051),
            .I(N__23048));
    Odrv4 I__2895 (
            .O(N__23048),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__2894 (
            .O(N__23045),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__2893 (
            .O(N__23042),
            .I(N__23039));
    LocalMux I__2892 (
            .O(N__23039),
            .I(N__23036));
    Span4Mux_v I__2891 (
            .O(N__23036),
            .I(N__23033));
    Sp12to4 I__2890 (
            .O(N__23033),
            .I(N__23030));
    Span12Mux_h I__2889 (
            .O(N__23030),
            .I(N__23027));
    Span12Mux_h I__2888 (
            .O(N__23027),
            .I(N__23024));
    Odrv12 I__2887 (
            .O(N__23024),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    CascadeMux I__2886 (
            .O(N__23021),
            .I(N__23018));
    InMux I__2885 (
            .O(N__23018),
            .I(N__23015));
    LocalMux I__2884 (
            .O(N__23015),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__2883 (
            .O(N__23012),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    InMux I__2882 (
            .O(N__23009),
            .I(N__23006));
    LocalMux I__2881 (
            .O(N__23006),
            .I(N__23003));
    Span4Mux_v I__2880 (
            .O(N__23003),
            .I(N__23000));
    Sp12to4 I__2879 (
            .O(N__23000),
            .I(N__22997));
    Span12Mux_h I__2878 (
            .O(N__22997),
            .I(N__22994));
    Span12Mux_v I__2877 (
            .O(N__22994),
            .I(N__22991));
    Odrv12 I__2876 (
            .O(N__22991),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__2875 (
            .O(N__22988),
            .I(N__22985));
    LocalMux I__2874 (
            .O(N__22985),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__2873 (
            .O(N__22982),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    CascadeMux I__2872 (
            .O(N__22979),
            .I(N__22976));
    InMux I__2871 (
            .O(N__22976),
            .I(N__22973));
    LocalMux I__2870 (
            .O(N__22973),
            .I(N__22970));
    Span4Mux_v I__2869 (
            .O(N__22970),
            .I(N__22967));
    Sp12to4 I__2868 (
            .O(N__22967),
            .I(N__22964));
    Span12Mux_h I__2867 (
            .O(N__22964),
            .I(N__22961));
    Span12Mux_h I__2866 (
            .O(N__22961),
            .I(N__22958));
    Odrv12 I__2865 (
            .O(N__22958),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    CascadeMux I__2864 (
            .O(N__22955),
            .I(N__22952));
    InMux I__2863 (
            .O(N__22952),
            .I(N__22949));
    LocalMux I__2862 (
            .O(N__22949),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__2861 (
            .O(N__22946),
            .I(bfn_5_15_0_));
    InMux I__2860 (
            .O(N__22943),
            .I(N__22940));
    LocalMux I__2859 (
            .O(N__22940),
            .I(N__22937));
    Span4Mux_h I__2858 (
            .O(N__22937),
            .I(N__22934));
    Sp12to4 I__2857 (
            .O(N__22934),
            .I(N__22931));
    Span12Mux_v I__2856 (
            .O(N__22931),
            .I(N__22928));
    Span12Mux_h I__2855 (
            .O(N__22928),
            .I(N__22925));
    Odrv12 I__2854 (
            .O(N__22925),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    CascadeMux I__2853 (
            .O(N__22922),
            .I(N__22919));
    InMux I__2852 (
            .O(N__22919),
            .I(N__22916));
    LocalMux I__2851 (
            .O(N__22916),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__2850 (
            .O(N__22913),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    CascadeMux I__2849 (
            .O(N__22910),
            .I(N__22907));
    InMux I__2848 (
            .O(N__22907),
            .I(N__22904));
    LocalMux I__2847 (
            .O(N__22904),
            .I(N__22901));
    Span4Mux_v I__2846 (
            .O(N__22901),
            .I(N__22898));
    Sp12to4 I__2845 (
            .O(N__22898),
            .I(N__22895));
    Span12Mux_h I__2844 (
            .O(N__22895),
            .I(N__22892));
    Span12Mux_h I__2843 (
            .O(N__22892),
            .I(N__22889));
    Odrv12 I__2842 (
            .O(N__22889),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__2841 (
            .O(N__22886),
            .I(N__22883));
    LocalMux I__2840 (
            .O(N__22883),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__2839 (
            .O(N__22880),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__2838 (
            .O(N__22877),
            .I(N__22874));
    LocalMux I__2837 (
            .O(N__22874),
            .I(N__22871));
    Span12Mux_h I__2836 (
            .O(N__22871),
            .I(N__22868));
    Span12Mux_h I__2835 (
            .O(N__22868),
            .I(N__22865));
    Odrv12 I__2834 (
            .O(N__22865),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    CascadeMux I__2833 (
            .O(N__22862),
            .I(N__22859));
    InMux I__2832 (
            .O(N__22859),
            .I(N__22856));
    LocalMux I__2831 (
            .O(N__22856),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__2830 (
            .O(N__22853),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__2829 (
            .O(N__22850),
            .I(N__22847));
    LocalMux I__2828 (
            .O(N__22847),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__2827 (
            .O(N__22844),
            .I(N__22841));
    LocalMux I__2826 (
            .O(N__22841),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    CascadeMux I__2825 (
            .O(N__22838),
            .I(N__22835));
    InMux I__2824 (
            .O(N__22835),
            .I(N__22832));
    LocalMux I__2823 (
            .O(N__22832),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__2822 (
            .O(N__22829),
            .I(N__22826));
    LocalMux I__2821 (
            .O(N__22826),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__2820 (
            .O(N__22823),
            .I(N__22820));
    LocalMux I__2819 (
            .O(N__22820),
            .I(N__22817));
    Span4Mux_h I__2818 (
            .O(N__22817),
            .I(N__22814));
    Span4Mux_h I__2817 (
            .O(N__22814),
            .I(N__22811));
    Odrv4 I__2816 (
            .O(N__22811),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    CascadeMux I__2815 (
            .O(N__22808),
            .I(N__22805));
    InMux I__2814 (
            .O(N__22805),
            .I(N__22802));
    LocalMux I__2813 (
            .O(N__22802),
            .I(N__22799));
    Span4Mux_v I__2812 (
            .O(N__22799),
            .I(N__22796));
    Sp12to4 I__2811 (
            .O(N__22796),
            .I(N__22793));
    Span12Mux_h I__2810 (
            .O(N__22793),
            .I(N__22790));
    Span12Mux_h I__2809 (
            .O(N__22790),
            .I(N__22787));
    Odrv12 I__2808 (
            .O(N__22787),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__2807 (
            .O(N__22784),
            .I(N__22781));
    InMux I__2806 (
            .O(N__22781),
            .I(N__22778));
    LocalMux I__2805 (
            .O(N__22778),
            .I(N__22775));
    Odrv4 I__2804 (
            .O(N__22775),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__2803 (
            .O(N__22772),
            .I(N__22769));
    LocalMux I__2802 (
            .O(N__22769),
            .I(N__22766));
    Span4Mux_h I__2801 (
            .O(N__22766),
            .I(N__22763));
    Sp12to4 I__2800 (
            .O(N__22763),
            .I(N__22760));
    Span12Mux_v I__2799 (
            .O(N__22760),
            .I(N__22757));
    Span12Mux_h I__2798 (
            .O(N__22757),
            .I(N__22754));
    Odrv12 I__2797 (
            .O(N__22754),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__2796 (
            .O(N__22751),
            .I(N__22748));
    InMux I__2795 (
            .O(N__22748),
            .I(N__22745));
    LocalMux I__2794 (
            .O(N__22745),
            .I(N__22742));
    Span4Mux_h I__2793 (
            .O(N__22742),
            .I(N__22739));
    Span4Mux_h I__2792 (
            .O(N__22739),
            .I(N__22736));
    Odrv4 I__2791 (
            .O(N__22736),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    CascadeMux I__2790 (
            .O(N__22733),
            .I(N__22730));
    InMux I__2789 (
            .O(N__22730),
            .I(N__22727));
    LocalMux I__2788 (
            .O(N__22727),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__2787 (
            .O(N__22724),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__2786 (
            .O(N__22721),
            .I(N__22718));
    LocalMux I__2785 (
            .O(N__22718),
            .I(N__22715));
    Span4Mux_v I__2784 (
            .O(N__22715),
            .I(N__22712));
    Sp12to4 I__2783 (
            .O(N__22712),
            .I(N__22709));
    Span12Mux_h I__2782 (
            .O(N__22709),
            .I(N__22706));
    Span12Mux_v I__2781 (
            .O(N__22706),
            .I(N__22703));
    Odrv12 I__2780 (
            .O(N__22703),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__2779 (
            .O(N__22700),
            .I(N__22697));
    InMux I__2778 (
            .O(N__22697),
            .I(N__22694));
    LocalMux I__2777 (
            .O(N__22694),
            .I(N__22691));
    Span4Mux_h I__2776 (
            .O(N__22691),
            .I(N__22688));
    Span4Mux_h I__2775 (
            .O(N__22688),
            .I(N__22685));
    Odrv4 I__2774 (
            .O(N__22685),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    CascadeMux I__2773 (
            .O(N__22682),
            .I(N__22679));
    InMux I__2772 (
            .O(N__22679),
            .I(N__22676));
    LocalMux I__2771 (
            .O(N__22676),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__2770 (
            .O(N__22673),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    InMux I__2769 (
            .O(N__22670),
            .I(N__22667));
    LocalMux I__2768 (
            .O(N__22667),
            .I(N__22664));
    Span12Mux_h I__2767 (
            .O(N__22664),
            .I(N__22661));
    Span12Mux_v I__2766 (
            .O(N__22661),
            .I(N__22658));
    Span12Mux_h I__2765 (
            .O(N__22658),
            .I(N__22655));
    Odrv12 I__2764 (
            .O(N__22655),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__2763 (
            .O(N__22652),
            .I(N__22649));
    InMux I__2762 (
            .O(N__22649),
            .I(N__22646));
    LocalMux I__2761 (
            .O(N__22646),
            .I(N__22643));
    Span12Mux_h I__2760 (
            .O(N__22643),
            .I(N__22640));
    Odrv12 I__2759 (
            .O(N__22640),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__2758 (
            .O(N__22637),
            .I(N__22634));
    LocalMux I__2757 (
            .O(N__22634),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__2756 (
            .O(N__22631),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    CascadeMux I__2755 (
            .O(N__22628),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__2754 (
            .O(N__22625),
            .I(N__22622));
    LocalMux I__2753 (
            .O(N__22622),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2752 (
            .O(N__22619),
            .I(N__22616));
    LocalMux I__2751 (
            .O(N__22616),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__2750 (
            .O(N__22613),
            .I(N__22610));
    LocalMux I__2749 (
            .O(N__22610),
            .I(N__22607));
    Odrv4 I__2748 (
            .O(N__22607),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__2747 (
            .O(N__22604),
            .I(N__22601));
    LocalMux I__2746 (
            .O(N__22601),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    CascadeMux I__2745 (
            .O(N__22598),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ));
    InMux I__2744 (
            .O(N__22595),
            .I(N__22592));
    LocalMux I__2743 (
            .O(N__22592),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2742 (
            .O(N__22589),
            .I(N__22585));
    InMux I__2741 (
            .O(N__22588),
            .I(N__22582));
    LocalMux I__2740 (
            .O(N__22585),
            .I(N__22579));
    LocalMux I__2739 (
            .O(N__22582),
            .I(N__22576));
    Span4Mux_h I__2738 (
            .O(N__22579),
            .I(N__22573));
    Odrv4 I__2737 (
            .O(N__22576),
            .I(pwm_duty_input_0));
    Odrv4 I__2736 (
            .O(N__22573),
            .I(pwm_duty_input_0));
    InMux I__2735 (
            .O(N__22568),
            .I(N__22565));
    LocalMux I__2734 (
            .O(N__22565),
            .I(N__22562));
    Odrv12 I__2733 (
            .O(N__22562),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2732 (
            .O(N__22559),
            .I(N__22555));
    InMux I__2731 (
            .O(N__22558),
            .I(N__22552));
    LocalMux I__2730 (
            .O(N__22555),
            .I(N__22549));
    LocalMux I__2729 (
            .O(N__22552),
            .I(N__22546));
    Span4Mux_h I__2728 (
            .O(N__22549),
            .I(N__22543));
    Odrv4 I__2727 (
            .O(N__22546),
            .I(pwm_duty_input_1));
    Odrv4 I__2726 (
            .O(N__22543),
            .I(pwm_duty_input_1));
    InMux I__2725 (
            .O(N__22538),
            .I(N__22535));
    LocalMux I__2724 (
            .O(N__22535),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__2723 (
            .O(N__22532),
            .I(N__22529));
    LocalMux I__2722 (
            .O(N__22529),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    CascadeMux I__2721 (
            .O(N__22526),
            .I(N__22523));
    InMux I__2720 (
            .O(N__22523),
            .I(N__22520));
    LocalMux I__2719 (
            .O(N__22520),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__2718 (
            .O(N__22517),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__2717 (
            .O(N__22514),
            .I(N__22511));
    LocalMux I__2716 (
            .O(N__22511),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__2715 (
            .O(N__22508),
            .I(N__22505));
    LocalMux I__2714 (
            .O(N__22505),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__2713 (
            .O(N__22502),
            .I(N__22499));
    InMux I__2712 (
            .O(N__22499),
            .I(N__22496));
    LocalMux I__2711 (
            .O(N__22496),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__2710 (
            .O(N__22493),
            .I(N__22490));
    LocalMux I__2709 (
            .O(N__22490),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__2708 (
            .O(N__22487),
            .I(N__22484));
    LocalMux I__2707 (
            .O(N__22484),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    CascadeMux I__2706 (
            .O(N__22481),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ));
    InMux I__2705 (
            .O(N__22478),
            .I(N__22475));
    LocalMux I__2704 (
            .O(N__22475),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    InMux I__2703 (
            .O(N__22472),
            .I(N__22469));
    LocalMux I__2702 (
            .O(N__22469),
            .I(\current_shift_inst.PI_CTRL.N_77 ));
    InMux I__2701 (
            .O(N__22466),
            .I(N__22463));
    LocalMux I__2700 (
            .O(N__22463),
            .I(N__22460));
    Odrv4 I__2699 (
            .O(N__22460),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    CascadeMux I__2698 (
            .O(N__22457),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ));
    CascadeMux I__2697 (
            .O(N__22454),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ));
    InMux I__2696 (
            .O(N__22451),
            .I(N__22448));
    LocalMux I__2695 (
            .O(N__22448),
            .I(N__22445));
    Odrv4 I__2694 (
            .O(N__22445),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    CascadeMux I__2693 (
            .O(N__22442),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__2692 (
            .O(N__22439),
            .I(N__22436));
    LocalMux I__2691 (
            .O(N__22436),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    CascadeMux I__2690 (
            .O(N__22433),
            .I(N__22430));
    InMux I__2689 (
            .O(N__22430),
            .I(N__22427));
    LocalMux I__2688 (
            .O(N__22427),
            .I(N__22424));
    Odrv12 I__2687 (
            .O(N__22424),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__2686 (
            .O(N__22421),
            .I(N__22418));
    LocalMux I__2685 (
            .O(N__22418),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    CascadeMux I__2684 (
            .O(N__22415),
            .I(N__22412));
    InMux I__2683 (
            .O(N__22412),
            .I(N__22409));
    LocalMux I__2682 (
            .O(N__22409),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__2681 (
            .O(N__22406),
            .I(N__22403));
    LocalMux I__2680 (
            .O(N__22403),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__2679 (
            .O(N__22400),
            .I(N__22397));
    LocalMux I__2678 (
            .O(N__22397),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    CascadeMux I__2677 (
            .O(N__22394),
            .I(N__22391));
    InMux I__2676 (
            .O(N__22391),
            .I(N__22388));
    LocalMux I__2675 (
            .O(N__22388),
            .I(N__22385));
    Span4Mux_h I__2674 (
            .O(N__22385),
            .I(N__22382));
    Odrv4 I__2673 (
            .O(N__22382),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__2672 (
            .O(N__22379),
            .I(N__22376));
    LocalMux I__2671 (
            .O(N__22376),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    CascadeMux I__2670 (
            .O(N__22373),
            .I(N__22370));
    InMux I__2669 (
            .O(N__22370),
            .I(N__22367));
    LocalMux I__2668 (
            .O(N__22367),
            .I(N__22364));
    Span4Mux_h I__2667 (
            .O(N__22364),
            .I(N__22361));
    Odrv4 I__2666 (
            .O(N__22361),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ));
    InMux I__2665 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__2664 (
            .O(N__22355),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    InMux I__2663 (
            .O(N__22352),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    InMux I__2662 (
            .O(N__22349),
            .I(bfn_4_15_0_));
    InMux I__2661 (
            .O(N__22346),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    InMux I__2660 (
            .O(N__22343),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    InMux I__2659 (
            .O(N__22340),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    InMux I__2658 (
            .O(N__22337),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    InMux I__2657 (
            .O(N__22334),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__2656 (
            .O(N__22331),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    CascadeMux I__2655 (
            .O(N__22328),
            .I(N__22325));
    InMux I__2654 (
            .O(N__22325),
            .I(N__22322));
    LocalMux I__2653 (
            .O(N__22322),
            .I(N__22319));
    Odrv4 I__2652 (
            .O(N__22319),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__2651 (
            .O(N__22316),
            .I(N__22313));
    InMux I__2650 (
            .O(N__22313),
            .I(N__22310));
    LocalMux I__2649 (
            .O(N__22310),
            .I(N__22307));
    Odrv4 I__2648 (
            .O(N__22307),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__2647 (
            .O(N__22304),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    InMux I__2646 (
            .O(N__22301),
            .I(bfn_4_14_0_));
    InMux I__2645 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__2644 (
            .O(N__22295),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__2643 (
            .O(N__22292),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__2642 (
            .O(N__22289),
            .I(N__22286));
    InMux I__2641 (
            .O(N__22286),
            .I(N__22283));
    LocalMux I__2640 (
            .O(N__22283),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__2639 (
            .O(N__22280),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__2638 (
            .O(N__22277),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    InMux I__2637 (
            .O(N__22274),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    InMux I__2636 (
            .O(N__22271),
            .I(N__22268));
    LocalMux I__2635 (
            .O(N__22268),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__2634 (
            .O(N__22265),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__2633 (
            .O(N__22262),
            .I(N__22259));
    InMux I__2632 (
            .O(N__22259),
            .I(N__22256));
    LocalMux I__2631 (
            .O(N__22256),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__2630 (
            .O(N__22253),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__2629 (
            .O(N__22250),
            .I(N__22247));
    InMux I__2628 (
            .O(N__22247),
            .I(N__22244));
    LocalMux I__2627 (
            .O(N__22244),
            .I(N__22241));
    Span4Mux_h I__2626 (
            .O(N__22241),
            .I(N__22238));
    Span4Mux_h I__2625 (
            .O(N__22238),
            .I(N__22235));
    Odrv4 I__2624 (
            .O(N__22235),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__2623 (
            .O(N__22232),
            .I(N__22229));
    LocalMux I__2622 (
            .O(N__22229),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__2621 (
            .O(N__22226),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    CascadeMux I__2620 (
            .O(N__22223),
            .I(N__22220));
    InMux I__2619 (
            .O(N__22220),
            .I(N__22217));
    LocalMux I__2618 (
            .O(N__22217),
            .I(N__22214));
    Span4Mux_v I__2617 (
            .O(N__22214),
            .I(N__22211));
    Odrv4 I__2616 (
            .O(N__22211),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    CascadeMux I__2615 (
            .O(N__22208),
            .I(N__22205));
    InMux I__2614 (
            .O(N__22205),
            .I(N__22202));
    LocalMux I__2613 (
            .O(N__22202),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__2612 (
            .O(N__22199),
            .I(bfn_4_13_0_));
    CascadeMux I__2611 (
            .O(N__22196),
            .I(N__22193));
    InMux I__2610 (
            .O(N__22193),
            .I(N__22190));
    LocalMux I__2609 (
            .O(N__22190),
            .I(N__22187));
    Span4Mux_v I__2608 (
            .O(N__22187),
            .I(N__22184));
    Odrv4 I__2607 (
            .O(N__22184),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__2606 (
            .O(N__22181),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__2605 (
            .O(N__22178),
            .I(N__22175));
    InMux I__2604 (
            .O(N__22175),
            .I(N__22172));
    LocalMux I__2603 (
            .O(N__22172),
            .I(N__22169));
    Span4Mux_v I__2602 (
            .O(N__22169),
            .I(N__22166));
    Span4Mux_h I__2601 (
            .O(N__22166),
            .I(N__22163));
    Odrv4 I__2600 (
            .O(N__22163),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    CascadeMux I__2599 (
            .O(N__22160),
            .I(N__22157));
    InMux I__2598 (
            .O(N__22157),
            .I(N__22154));
    LocalMux I__2597 (
            .O(N__22154),
            .I(N__22151));
    Span4Mux_h I__2596 (
            .O(N__22151),
            .I(N__22148));
    Odrv4 I__2595 (
            .O(N__22148),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__2594 (
            .O(N__22145),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__2593 (
            .O(N__22142),
            .I(N__22139));
    LocalMux I__2592 (
            .O(N__22139),
            .I(N__22136));
    Span4Mux_v I__2591 (
            .O(N__22136),
            .I(N__22133));
    Odrv4 I__2590 (
            .O(N__22133),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__2589 (
            .O(N__22130),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__2588 (
            .O(N__22127),
            .I(N__22124));
    InMux I__2587 (
            .O(N__22124),
            .I(N__22121));
    LocalMux I__2586 (
            .O(N__22121),
            .I(N__22118));
    Span4Mux_v I__2585 (
            .O(N__22118),
            .I(N__22115));
    Odrv4 I__2584 (
            .O(N__22115),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__2583 (
            .O(N__22112),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    CascadeMux I__2582 (
            .O(N__22109),
            .I(N__22106));
    InMux I__2581 (
            .O(N__22106),
            .I(N__22103));
    LocalMux I__2580 (
            .O(N__22103),
            .I(N__22100));
    Span4Mux_h I__2579 (
            .O(N__22100),
            .I(N__22097));
    Odrv4 I__2578 (
            .O(N__22097),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__2577 (
            .O(N__22094),
            .I(N__22091));
    LocalMux I__2576 (
            .O(N__22091),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__2575 (
            .O(N__22088),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    InMux I__2574 (
            .O(N__22085),
            .I(N__22082));
    LocalMux I__2573 (
            .O(N__22082),
            .I(N__22079));
    Span4Mux_h I__2572 (
            .O(N__22079),
            .I(N__22076));
    Odrv4 I__2571 (
            .O(N__22076),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    CascadeMux I__2570 (
            .O(N__22073),
            .I(N__22070));
    InMux I__2569 (
            .O(N__22070),
            .I(N__22067));
    LocalMux I__2568 (
            .O(N__22067),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__2567 (
            .O(N__22064),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    InMux I__2566 (
            .O(N__22061),
            .I(N__22058));
    LocalMux I__2565 (
            .O(N__22058),
            .I(N__22053));
    InMux I__2564 (
            .O(N__22057),
            .I(N__22048));
    InMux I__2563 (
            .O(N__22056),
            .I(N__22048));
    Span4Mux_s3_h I__2562 (
            .O(N__22053),
            .I(N__22045));
    LocalMux I__2561 (
            .O(N__22048),
            .I(pwm_duty_input_7));
    Odrv4 I__2560 (
            .O(N__22045),
            .I(pwm_duty_input_7));
    CascadeMux I__2559 (
            .O(N__22040),
            .I(N__22036));
    InMux I__2558 (
            .O(N__22039),
            .I(N__22033));
    InMux I__2557 (
            .O(N__22036),
            .I(N__22030));
    LocalMux I__2556 (
            .O(N__22033),
            .I(N__22025));
    LocalMux I__2555 (
            .O(N__22030),
            .I(N__22025));
    Span4Mux_v I__2554 (
            .O(N__22025),
            .I(N__22022));
    Odrv4 I__2553 (
            .O(N__22022),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    InMux I__2552 (
            .O(N__22019),
            .I(N__22016));
    LocalMux I__2551 (
            .O(N__22016),
            .I(N__22013));
    Span4Mux_v I__2550 (
            .O(N__22013),
            .I(N__22010));
    Odrv4 I__2549 (
            .O(N__22010),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__2548 (
            .O(N__22007),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    CascadeMux I__2547 (
            .O(N__22004),
            .I(N__22001));
    InMux I__2546 (
            .O(N__22001),
            .I(N__21998));
    LocalMux I__2545 (
            .O(N__21998),
            .I(N__21995));
    Span4Mux_v I__2544 (
            .O(N__21995),
            .I(N__21992));
    Odrv4 I__2543 (
            .O(N__21992),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__2542 (
            .O(N__21989),
            .I(N__21986));
    LocalMux I__2541 (
            .O(N__21986),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__2540 (
            .O(N__21983),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    InMux I__2539 (
            .O(N__21980),
            .I(N__21977));
    LocalMux I__2538 (
            .O(N__21977),
            .I(N__21974));
    Span4Mux_v I__2537 (
            .O(N__21974),
            .I(N__21971));
    Odrv4 I__2536 (
            .O(N__21971),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    InMux I__2535 (
            .O(N__21968),
            .I(N__21965));
    LocalMux I__2534 (
            .O(N__21965),
            .I(N__21962));
    Span4Mux_h I__2533 (
            .O(N__21962),
            .I(N__21959));
    Odrv4 I__2532 (
            .O(N__21959),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__2531 (
            .O(N__21956),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__2530 (
            .O(N__21953),
            .I(N__21950));
    InMux I__2529 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__2528 (
            .O(N__21947),
            .I(N__21944));
    Span4Mux_v I__2527 (
            .O(N__21944),
            .I(N__21941));
    Odrv4 I__2526 (
            .O(N__21941),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    CascadeMux I__2525 (
            .O(N__21938),
            .I(N__21935));
    InMux I__2524 (
            .O(N__21935),
            .I(N__21932));
    LocalMux I__2523 (
            .O(N__21932),
            .I(N__21929));
    Span4Mux_v I__2522 (
            .O(N__21929),
            .I(N__21926));
    Odrv4 I__2521 (
            .O(N__21926),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__2520 (
            .O(N__21923),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__2519 (
            .O(N__21920),
            .I(N__21917));
    InMux I__2518 (
            .O(N__21917),
            .I(N__21914));
    LocalMux I__2517 (
            .O(N__21914),
            .I(N__21911));
    Span4Mux_v I__2516 (
            .O(N__21911),
            .I(N__21908));
    Odrv4 I__2515 (
            .O(N__21908),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__2514 (
            .O(N__21905),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__2513 (
            .O(N__21902),
            .I(N__21899));
    InMux I__2512 (
            .O(N__21899),
            .I(N__21896));
    LocalMux I__2511 (
            .O(N__21896),
            .I(N__21893));
    Span4Mux_h I__2510 (
            .O(N__21893),
            .I(N__21890));
    Odrv4 I__2509 (
            .O(N__21890),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__2508 (
            .O(N__21887),
            .I(N__21884));
    LocalMux I__2507 (
            .O(N__21884),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__2506 (
            .O(N__21881),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__2505 (
            .O(N__21878),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__2504 (
            .O(N__21875),
            .I(N__21872));
    LocalMux I__2503 (
            .O(N__21872),
            .I(N__21869));
    Odrv4 I__2502 (
            .O(N__21869),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    InMux I__2501 (
            .O(N__21866),
            .I(N__21863));
    LocalMux I__2500 (
            .O(N__21863),
            .I(N__21860));
    Odrv4 I__2499 (
            .O(N__21860),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    CascadeMux I__2498 (
            .O(N__21857),
            .I(\current_shift_inst.PI_CTRL.N_98_cascade_ ));
    InMux I__2497 (
            .O(N__21854),
            .I(N__21851));
    LocalMux I__2496 (
            .O(N__21851),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    CascadeMux I__2495 (
            .O(N__21848),
            .I(\current_shift_inst.PI_CTRL.N_96_cascade_ ));
    InMux I__2494 (
            .O(N__21845),
            .I(N__21841));
    CascadeMux I__2493 (
            .O(N__21844),
            .I(N__21838));
    LocalMux I__2492 (
            .O(N__21841),
            .I(N__21834));
    InMux I__2491 (
            .O(N__21838),
            .I(N__21829));
    InMux I__2490 (
            .O(N__21837),
            .I(N__21829));
    Span4Mux_s3_h I__2489 (
            .O(N__21834),
            .I(N__21826));
    LocalMux I__2488 (
            .O(N__21829),
            .I(pwm_duty_input_6));
    Odrv4 I__2487 (
            .O(N__21826),
            .I(pwm_duty_input_6));
    InMux I__2486 (
            .O(N__21821),
            .I(N__21818));
    LocalMux I__2485 (
            .O(N__21818),
            .I(N__21815));
    Odrv4 I__2484 (
            .O(N__21815),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__2483 (
            .O(N__21812),
            .I(N__21809));
    InMux I__2482 (
            .O(N__21809),
            .I(N__21805));
    InMux I__2481 (
            .O(N__21808),
            .I(N__21802));
    LocalMux I__2480 (
            .O(N__21805),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__2479 (
            .O(N__21802),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__2478 (
            .O(N__21797),
            .I(N__21794));
    InMux I__2477 (
            .O(N__21794),
            .I(N__21789));
    InMux I__2476 (
            .O(N__21793),
            .I(N__21786));
    InMux I__2475 (
            .O(N__21792),
            .I(N__21783));
    LocalMux I__2474 (
            .O(N__21789),
            .I(N__21780));
    LocalMux I__2473 (
            .O(N__21786),
            .I(N__21777));
    LocalMux I__2472 (
            .O(N__21783),
            .I(N__21774));
    Span4Mux_v I__2471 (
            .O(N__21780),
            .I(N__21767));
    Span4Mux_v I__2470 (
            .O(N__21777),
            .I(N__21767));
    Span4Mux_s3_h I__2469 (
            .O(N__21774),
            .I(N__21767));
    Odrv4 I__2468 (
            .O(N__21767),
            .I(pwm_duty_input_4));
    InMux I__2467 (
            .O(N__21764),
            .I(N__21760));
    InMux I__2466 (
            .O(N__21763),
            .I(N__21757));
    LocalMux I__2465 (
            .O(N__21760),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    LocalMux I__2464 (
            .O(N__21757),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    InMux I__2463 (
            .O(N__21752),
            .I(N__21749));
    LocalMux I__2462 (
            .O(N__21749),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__2461 (
            .O(N__21746),
            .I(N__21741));
    InMux I__2460 (
            .O(N__21745),
            .I(N__21738));
    InMux I__2459 (
            .O(N__21744),
            .I(N__21735));
    LocalMux I__2458 (
            .O(N__21741),
            .I(N__21732));
    LocalMux I__2457 (
            .O(N__21738),
            .I(N__21727));
    LocalMux I__2456 (
            .O(N__21735),
            .I(N__21727));
    Span4Mux_s3_h I__2455 (
            .O(N__21732),
            .I(N__21724));
    Odrv4 I__2454 (
            .O(N__21727),
            .I(pwm_duty_input_3));
    Odrv4 I__2453 (
            .O(N__21724),
            .I(pwm_duty_input_3));
    CascadeMux I__2452 (
            .O(N__21719),
            .I(N__21715));
    InMux I__2451 (
            .O(N__21718),
            .I(N__21712));
    InMux I__2450 (
            .O(N__21715),
            .I(N__21709));
    LocalMux I__2449 (
            .O(N__21712),
            .I(N__21705));
    LocalMux I__2448 (
            .O(N__21709),
            .I(N__21702));
    InMux I__2447 (
            .O(N__21708),
            .I(N__21699));
    Span4Mux_s3_h I__2446 (
            .O(N__21705),
            .I(N__21696));
    Odrv12 I__2445 (
            .O(N__21702),
            .I(pwm_duty_input_5));
    LocalMux I__2444 (
            .O(N__21699),
            .I(pwm_duty_input_5));
    Odrv4 I__2443 (
            .O(N__21696),
            .I(pwm_duty_input_5));
    CascadeMux I__2442 (
            .O(N__21689),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11_cascade_ ));
    CascadeMux I__2441 (
            .O(N__21686),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    CascadeMux I__2440 (
            .O(N__21683),
            .I(\current_shift_inst.PI_CTRL.N_31_cascade_ ));
    InMux I__2439 (
            .O(N__21680),
            .I(N__21677));
    LocalMux I__2438 (
            .O(N__21677),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ));
    InMux I__2437 (
            .O(N__21674),
            .I(N__21670));
    InMux I__2436 (
            .O(N__21673),
            .I(N__21667));
    LocalMux I__2435 (
            .O(N__21670),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__2434 (
            .O(N__21667),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__2433 (
            .O(N__21662),
            .I(N__21659));
    InMux I__2432 (
            .O(N__21659),
            .I(N__21656));
    LocalMux I__2431 (
            .O(N__21656),
            .I(\pwm_generator_inst.threshold_9 ));
    InMux I__2430 (
            .O(N__21653),
            .I(N__21650));
    LocalMux I__2429 (
            .O(N__21650),
            .I(N__21646));
    InMux I__2428 (
            .O(N__21649),
            .I(N__21642));
    Span4Mux_h I__2427 (
            .O(N__21646),
            .I(N__21639));
    InMux I__2426 (
            .O(N__21645),
            .I(N__21636));
    LocalMux I__2425 (
            .O(N__21642),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__2424 (
            .O(N__21639),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2423 (
            .O(N__21636),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__2422 (
            .O(N__21629),
            .I(N__21626));
    LocalMux I__2421 (
            .O(N__21626),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2420 (
            .O(N__21623),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2419 (
            .O(N__21620),
            .I(N__21617));
    LocalMux I__2418 (
            .O(N__21617),
            .I(N__21614));
    Span4Mux_s2_v I__2417 (
            .O(N__21614),
            .I(N__21611));
    Sp12to4 I__2416 (
            .O(N__21611),
            .I(N__21608));
    Span12Mux_s10_h I__2415 (
            .O(N__21608),
            .I(N__21605));
    Span12Mux_h I__2414 (
            .O(N__21605),
            .I(N__21602));
    Span12Mux_v I__2413 (
            .O(N__21602),
            .I(N__21599));
    Odrv12 I__2412 (
            .O(N__21599),
            .I(pwm_output_c));
    CascadeMux I__2411 (
            .O(N__21596),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__2410 (
            .O(N__21593),
            .I(N__21573));
    InMux I__2409 (
            .O(N__21592),
            .I(N__21573));
    InMux I__2408 (
            .O(N__21591),
            .I(N__21573));
    InMux I__2407 (
            .O(N__21590),
            .I(N__21573));
    InMux I__2406 (
            .O(N__21589),
            .I(N__21573));
    InMux I__2405 (
            .O(N__21588),
            .I(N__21564));
    InMux I__2404 (
            .O(N__21587),
            .I(N__21564));
    InMux I__2403 (
            .O(N__21586),
            .I(N__21564));
    InMux I__2402 (
            .O(N__21585),
            .I(N__21564));
    InMux I__2401 (
            .O(N__21584),
            .I(N__21561));
    LocalMux I__2400 (
            .O(N__21573),
            .I(N__21558));
    LocalMux I__2399 (
            .O(N__21564),
            .I(N__21555));
    LocalMux I__2398 (
            .O(N__21561),
            .I(N__21548));
    Span4Mux_v I__2397 (
            .O(N__21558),
            .I(N__21548));
    Span4Mux_s3_h I__2396 (
            .O(N__21555),
            .I(N__21548));
    Odrv4 I__2395 (
            .O(N__21548),
            .I(\pwm_generator_inst.N_17 ));
    InMux I__2394 (
            .O(N__21545),
            .I(N__21542));
    LocalMux I__2393 (
            .O(N__21542),
            .I(N__21539));
    Odrv4 I__2392 (
            .O(N__21539),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__2391 (
            .O(N__21536),
            .I(N__21533));
    InMux I__2390 (
            .O(N__21533),
            .I(N__21530));
    LocalMux I__2389 (
            .O(N__21530),
            .I(N__21527));
    Odrv4 I__2388 (
            .O(N__21527),
            .I(\pwm_generator_inst.threshold_2 ));
    InMux I__2387 (
            .O(N__21524),
            .I(N__21521));
    LocalMux I__2386 (
            .O(N__21521),
            .I(N__21517));
    InMux I__2385 (
            .O(N__21520),
            .I(N__21513));
    Span4Mux_h I__2384 (
            .O(N__21517),
            .I(N__21510));
    InMux I__2383 (
            .O(N__21516),
            .I(N__21507));
    LocalMux I__2382 (
            .O(N__21513),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__2381 (
            .O(N__21510),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2380 (
            .O(N__21507),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2379 (
            .O(N__21500),
            .I(N__21497));
    LocalMux I__2378 (
            .O(N__21497),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__2377 (
            .O(N__21494),
            .I(N__21490));
    InMux I__2376 (
            .O(N__21493),
            .I(N__21486));
    LocalMux I__2375 (
            .O(N__21490),
            .I(N__21483));
    InMux I__2374 (
            .O(N__21489),
            .I(N__21480));
    LocalMux I__2373 (
            .O(N__21486),
            .I(N__21475));
    Span4Mux_v I__2372 (
            .O(N__21483),
            .I(N__21475));
    LocalMux I__2371 (
            .O(N__21480),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__2370 (
            .O(N__21475),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    CascadeMux I__2369 (
            .O(N__21470),
            .I(N__21467));
    InMux I__2368 (
            .O(N__21467),
            .I(N__21464));
    LocalMux I__2367 (
            .O(N__21464),
            .I(N__21461));
    Odrv12 I__2366 (
            .O(N__21461),
            .I(\pwm_generator_inst.threshold_3 ));
    InMux I__2365 (
            .O(N__21458),
            .I(N__21455));
    LocalMux I__2364 (
            .O(N__21455),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__2363 (
            .O(N__21452),
            .I(N__21449));
    LocalMux I__2362 (
            .O(N__21449),
            .I(N__21444));
    InMux I__2361 (
            .O(N__21448),
            .I(N__21441));
    InMux I__2360 (
            .O(N__21447),
            .I(N__21438));
    Span4Mux_v I__2359 (
            .O(N__21444),
            .I(N__21435));
    LocalMux I__2358 (
            .O(N__21441),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2357 (
            .O(N__21438),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__2356 (
            .O(N__21435),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    CascadeMux I__2355 (
            .O(N__21428),
            .I(N__21425));
    InMux I__2354 (
            .O(N__21425),
            .I(N__21422));
    LocalMux I__2353 (
            .O(N__21422),
            .I(\pwm_generator_inst.threshold_4 ));
    InMux I__2352 (
            .O(N__21419),
            .I(N__21416));
    LocalMux I__2351 (
            .O(N__21416),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__2350 (
            .O(N__21413),
            .I(N__21410));
    InMux I__2349 (
            .O(N__21410),
            .I(N__21407));
    LocalMux I__2348 (
            .O(N__21407),
            .I(N__21404));
    Odrv4 I__2347 (
            .O(N__21404),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__2346 (
            .O(N__21401),
            .I(N__21398));
    LocalMux I__2345 (
            .O(N__21398),
            .I(N__21393));
    InMux I__2344 (
            .O(N__21397),
            .I(N__21390));
    InMux I__2343 (
            .O(N__21396),
            .I(N__21387));
    Span4Mux_v I__2342 (
            .O(N__21393),
            .I(N__21384));
    LocalMux I__2341 (
            .O(N__21390),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2340 (
            .O(N__21387),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__2339 (
            .O(N__21384),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2338 (
            .O(N__21377),
            .I(N__21374));
    LocalMux I__2337 (
            .O(N__21374),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__2336 (
            .O(N__21371),
            .I(N__21368));
    InMux I__2335 (
            .O(N__21368),
            .I(N__21365));
    LocalMux I__2334 (
            .O(N__21365),
            .I(\pwm_generator_inst.un14_counter_6 ));
    InMux I__2333 (
            .O(N__21362),
            .I(N__21359));
    LocalMux I__2332 (
            .O(N__21359),
            .I(N__21354));
    InMux I__2331 (
            .O(N__21358),
            .I(N__21351));
    InMux I__2330 (
            .O(N__21357),
            .I(N__21348));
    Span4Mux_h I__2329 (
            .O(N__21354),
            .I(N__21345));
    LocalMux I__2328 (
            .O(N__21351),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2327 (
            .O(N__21348),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__2326 (
            .O(N__21345),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__2325 (
            .O(N__21338),
            .I(N__21335));
    LocalMux I__2324 (
            .O(N__21335),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2323 (
            .O(N__21332),
            .I(N__21329));
    InMux I__2322 (
            .O(N__21329),
            .I(N__21326));
    LocalMux I__2321 (
            .O(N__21326),
            .I(\pwm_generator_inst.un14_counter_7 ));
    InMux I__2320 (
            .O(N__21323),
            .I(N__21320));
    LocalMux I__2319 (
            .O(N__21320),
            .I(N__21315));
    InMux I__2318 (
            .O(N__21319),
            .I(N__21312));
    InMux I__2317 (
            .O(N__21318),
            .I(N__21309));
    Span4Mux_v I__2316 (
            .O(N__21315),
            .I(N__21306));
    LocalMux I__2315 (
            .O(N__21312),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2314 (
            .O(N__21309),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2313 (
            .O(N__21306),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2312 (
            .O(N__21299),
            .I(N__21296));
    LocalMux I__2311 (
            .O(N__21296),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2310 (
            .O(N__21293),
            .I(N__21290));
    InMux I__2309 (
            .O(N__21290),
            .I(N__21287));
    LocalMux I__2308 (
            .O(N__21287),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__2307 (
            .O(N__21284),
            .I(N__21281));
    LocalMux I__2306 (
            .O(N__21281),
            .I(N__21277));
    InMux I__2305 (
            .O(N__21280),
            .I(N__21273));
    Span4Mux_h I__2304 (
            .O(N__21277),
            .I(N__21270));
    InMux I__2303 (
            .O(N__21276),
            .I(N__21267));
    LocalMux I__2302 (
            .O(N__21273),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__2301 (
            .O(N__21270),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2300 (
            .O(N__21267),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2299 (
            .O(N__21260),
            .I(N__21257));
    LocalMux I__2298 (
            .O(N__21257),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__2297 (
            .O(N__21254),
            .I(N__21251));
    InMux I__2296 (
            .O(N__21251),
            .I(N__21248));
    LocalMux I__2295 (
            .O(N__21248),
            .I(N__21245));
    Odrv4 I__2294 (
            .O(N__21245),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__2293 (
            .O(N__21242),
            .I(N__21239));
    LocalMux I__2292 (
            .O(N__21239),
            .I(N__21235));
    InMux I__2291 (
            .O(N__21238),
            .I(N__21231));
    Span4Mux_h I__2290 (
            .O(N__21235),
            .I(N__21228));
    InMux I__2289 (
            .O(N__21234),
            .I(N__21225));
    LocalMux I__2288 (
            .O(N__21231),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__2287 (
            .O(N__21228),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2286 (
            .O(N__21225),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2285 (
            .O(N__21218),
            .I(N__21215));
    LocalMux I__2284 (
            .O(N__21215),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__2283 (
            .O(N__21212),
            .I(N__21209));
    InMux I__2282 (
            .O(N__21209),
            .I(N__21206));
    LocalMux I__2281 (
            .O(N__21206),
            .I(N__21203));
    Odrv4 I__2280 (
            .O(N__21203),
            .I(\pwm_generator_inst.un14_counter_1 ));
    InMux I__2279 (
            .O(N__21200),
            .I(N__21197));
    LocalMux I__2278 (
            .O(N__21197),
            .I(N__21192));
    InMux I__2277 (
            .O(N__21196),
            .I(N__21189));
    InMux I__2276 (
            .O(N__21195),
            .I(N__21186));
    Span4Mux_h I__2275 (
            .O(N__21192),
            .I(N__21183));
    LocalMux I__2274 (
            .O(N__21189),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2273 (
            .O(N__21186),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__2272 (
            .O(N__21183),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__2271 (
            .O(N__21176),
            .I(N__21172));
    InMux I__2270 (
            .O(N__21175),
            .I(N__21169));
    LocalMux I__2269 (
            .O(N__21172),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    LocalMux I__2268 (
            .O(N__21169),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    InMux I__2267 (
            .O(N__21164),
            .I(N__21161));
    LocalMux I__2266 (
            .O(N__21161),
            .I(N__21156));
    InMux I__2265 (
            .O(N__21160),
            .I(N__21151));
    InMux I__2264 (
            .O(N__21159),
            .I(N__21151));
    Odrv4 I__2263 (
            .O(N__21156),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__2262 (
            .O(N__21151),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    CascadeMux I__2261 (
            .O(N__21146),
            .I(N__21142));
    CascadeMux I__2260 (
            .O(N__21145),
            .I(N__21139));
    InMux I__2259 (
            .O(N__21142),
            .I(N__21136));
    InMux I__2258 (
            .O(N__21139),
            .I(N__21133));
    LocalMux I__2257 (
            .O(N__21136),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    LocalMux I__2256 (
            .O(N__21133),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    InMux I__2255 (
            .O(N__21128),
            .I(N__21125));
    LocalMux I__2254 (
            .O(N__21125),
            .I(N__21122));
    Span4Mux_s2_h I__2253 (
            .O(N__21122),
            .I(N__21117));
    InMux I__2252 (
            .O(N__21121),
            .I(N__21112));
    InMux I__2251 (
            .O(N__21120),
            .I(N__21112));
    Odrv4 I__2250 (
            .O(N__21117),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__2249 (
            .O(N__21112),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__2248 (
            .O(N__21107),
            .I(N__21104));
    LocalMux I__2247 (
            .O(N__21104),
            .I(N__21101));
    Odrv12 I__2246 (
            .O(N__21101),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__2245 (
            .O(N__21098),
            .I(N__21094));
    InMux I__2244 (
            .O(N__21097),
            .I(N__21091));
    LocalMux I__2243 (
            .O(N__21094),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    LocalMux I__2242 (
            .O(N__21091),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    InMux I__2241 (
            .O(N__21086),
            .I(N__21083));
    LocalMux I__2240 (
            .O(N__21083),
            .I(N__21078));
    InMux I__2239 (
            .O(N__21082),
            .I(N__21073));
    InMux I__2238 (
            .O(N__21081),
            .I(N__21073));
    Odrv4 I__2237 (
            .O(N__21078),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__2236 (
            .O(N__21073),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__2235 (
            .O(N__21068),
            .I(N__21065));
    LocalMux I__2234 (
            .O(N__21065),
            .I(N__21062));
    Odrv4 I__2233 (
            .O(N__21062),
            .I(un7_start_stop));
    CascadeMux I__2232 (
            .O(N__21059),
            .I(N__21056));
    InMux I__2231 (
            .O(N__21056),
            .I(N__21051));
    InMux I__2230 (
            .O(N__21055),
            .I(N__21048));
    InMux I__2229 (
            .O(N__21054),
            .I(N__21045));
    LocalMux I__2228 (
            .O(N__21051),
            .I(N__21042));
    LocalMux I__2227 (
            .O(N__21048),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__2226 (
            .O(N__21045),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv12 I__2225 (
            .O(N__21042),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__2224 (
            .O(N__21035),
            .I(N__21032));
    LocalMux I__2223 (
            .O(N__21032),
            .I(N__21029));
    Span4Mux_s3_h I__2222 (
            .O(N__21029),
            .I(N__21026));
    Odrv4 I__2221 (
            .O(N__21026),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__2220 (
            .O(N__21023),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__2219 (
            .O(N__21020),
            .I(N__21017));
    LocalMux I__2218 (
            .O(N__21017),
            .I(N__21012));
    InMux I__2217 (
            .O(N__21016),
            .I(N__21009));
    InMux I__2216 (
            .O(N__21015),
            .I(N__21006));
    Sp12to4 I__2215 (
            .O(N__21012),
            .I(N__21001));
    LocalMux I__2214 (
            .O(N__21009),
            .I(N__21001));
    LocalMux I__2213 (
            .O(N__21006),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    Odrv12 I__2212 (
            .O(N__21001),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    InMux I__2211 (
            .O(N__20996),
            .I(N__20993));
    LocalMux I__2210 (
            .O(N__20993),
            .I(N__20990));
    Span4Mux_s3_h I__2209 (
            .O(N__20990),
            .I(N__20987));
    Odrv4 I__2208 (
            .O(N__20987),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__2207 (
            .O(N__20984),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__2206 (
            .O(N__20981),
            .I(N__20978));
    LocalMux I__2205 (
            .O(N__20978),
            .I(N__20973));
    InMux I__2204 (
            .O(N__20977),
            .I(N__20970));
    InMux I__2203 (
            .O(N__20976),
            .I(N__20967));
    Span4Mux_v I__2202 (
            .O(N__20973),
            .I(N__20964));
    LocalMux I__2201 (
            .O(N__20970),
            .I(N__20961));
    LocalMux I__2200 (
            .O(N__20967),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__2199 (
            .O(N__20964),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__2198 (
            .O(N__20961),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__2197 (
            .O(N__20954),
            .I(N__20951));
    LocalMux I__2196 (
            .O(N__20951),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__2195 (
            .O(N__20948),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    CascadeMux I__2194 (
            .O(N__20945),
            .I(N__20940));
    InMux I__2193 (
            .O(N__20944),
            .I(N__20937));
    InMux I__2192 (
            .O(N__20943),
            .I(N__20934));
    InMux I__2191 (
            .O(N__20940),
            .I(N__20931));
    LocalMux I__2190 (
            .O(N__20937),
            .I(N__20928));
    LocalMux I__2189 (
            .O(N__20934),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__2188 (
            .O(N__20931),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv4 I__2187 (
            .O(N__20928),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__2186 (
            .O(N__20921),
            .I(N__20918));
    LocalMux I__2185 (
            .O(N__20918),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    InMux I__2184 (
            .O(N__20915),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__2183 (
            .O(N__20912),
            .I(N__20909));
    LocalMux I__2182 (
            .O(N__20909),
            .I(N__20906));
    Odrv4 I__2181 (
            .O(N__20906),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__2180 (
            .O(N__20903),
            .I(bfn_2_23_0_));
    CascadeMux I__2179 (
            .O(N__20900),
            .I(N__20897));
    InMux I__2178 (
            .O(N__20897),
            .I(N__20894));
    LocalMux I__2177 (
            .O(N__20894),
            .I(N__20891));
    Span4Mux_s2_h I__2176 (
            .O(N__20891),
            .I(N__20888));
    Odrv4 I__2175 (
            .O(N__20888),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__2174 (
            .O(N__20885),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__2173 (
            .O(N__20882),
            .I(N__20879));
    LocalMux I__2172 (
            .O(N__20879),
            .I(N__20876));
    Odrv4 I__2171 (
            .O(N__20876),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__2170 (
            .O(N__20873),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__2169 (
            .O(N__20870),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__2168 (
            .O(N__20867),
            .I(N__20864));
    LocalMux I__2167 (
            .O(N__20864),
            .I(N__20861));
    Span4Mux_v I__2166 (
            .O(N__20861),
            .I(N__20858));
    Odrv4 I__2165 (
            .O(N__20858),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__2164 (
            .O(N__20855),
            .I(N__20852));
    LocalMux I__2163 (
            .O(N__20852),
            .I(N__20849));
    Span4Mux_h I__2162 (
            .O(N__20849),
            .I(N__20846));
    Odrv4 I__2161 (
            .O(N__20846),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__2160 (
            .O(N__20843),
            .I(N__20840));
    LocalMux I__2159 (
            .O(N__20840),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__2158 (
            .O(N__20837),
            .I(N__20834));
    LocalMux I__2157 (
            .O(N__20834),
            .I(N__20831));
    Span4Mux_h I__2156 (
            .O(N__20831),
            .I(N__20828));
    Odrv4 I__2155 (
            .O(N__20828),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__2154 (
            .O(N__20825),
            .I(N__20822));
    LocalMux I__2153 (
            .O(N__20822),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__2152 (
            .O(N__20819),
            .I(N__20816));
    LocalMux I__2151 (
            .O(N__20816),
            .I(N__20813));
    Span4Mux_h I__2150 (
            .O(N__20813),
            .I(N__20810));
    Odrv4 I__2149 (
            .O(N__20810),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__2148 (
            .O(N__20807),
            .I(N__20804));
    LocalMux I__2147 (
            .O(N__20804),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__2146 (
            .O(N__20801),
            .I(N__20798));
    LocalMux I__2145 (
            .O(N__20798),
            .I(N__20795));
    Span4Mux_h I__2144 (
            .O(N__20795),
            .I(N__20792));
    Odrv4 I__2143 (
            .O(N__20792),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__2142 (
            .O(N__20789),
            .I(N__20786));
    LocalMux I__2141 (
            .O(N__20786),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__2140 (
            .O(N__20783),
            .I(N__20780));
    LocalMux I__2139 (
            .O(N__20780),
            .I(N__20777));
    Span4Mux_h I__2138 (
            .O(N__20777),
            .I(N__20774));
    Odrv4 I__2137 (
            .O(N__20774),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__2136 (
            .O(N__20771),
            .I(N__20768));
    LocalMux I__2135 (
            .O(N__20768),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__2134 (
            .O(N__20765),
            .I(N__20762));
    LocalMux I__2133 (
            .O(N__20762),
            .I(N__20759));
    Span4Mux_h I__2132 (
            .O(N__20759),
            .I(N__20756));
    Odrv4 I__2131 (
            .O(N__20756),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__2130 (
            .O(N__20753),
            .I(N__20750));
    LocalMux I__2129 (
            .O(N__20750),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__2128 (
            .O(N__20747),
            .I(N__20742));
    InMux I__2127 (
            .O(N__20746),
            .I(N__20739));
    InMux I__2126 (
            .O(N__20745),
            .I(N__20736));
    LocalMux I__2125 (
            .O(N__20742),
            .I(N__20733));
    LocalMux I__2124 (
            .O(N__20739),
            .I(N__20730));
    LocalMux I__2123 (
            .O(N__20736),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__2122 (
            .O(N__20733),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv12 I__2121 (
            .O(N__20730),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__2120 (
            .O(N__20723),
            .I(N__20720));
    LocalMux I__2119 (
            .O(N__20720),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    InMux I__2118 (
            .O(N__20717),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    CascadeMux I__2117 (
            .O(N__20714),
            .I(N__20710));
    CascadeMux I__2116 (
            .O(N__20713),
            .I(N__20704));
    InMux I__2115 (
            .O(N__20710),
            .I(N__20699));
    CascadeMux I__2114 (
            .O(N__20709),
            .I(N__20696));
    CascadeMux I__2113 (
            .O(N__20708),
            .I(N__20692));
    InMux I__2112 (
            .O(N__20707),
            .I(N__20686));
    InMux I__2111 (
            .O(N__20704),
            .I(N__20683));
    InMux I__2110 (
            .O(N__20703),
            .I(N__20678));
    InMux I__2109 (
            .O(N__20702),
            .I(N__20678));
    LocalMux I__2108 (
            .O(N__20699),
            .I(N__20675));
    InMux I__2107 (
            .O(N__20696),
            .I(N__20668));
    InMux I__2106 (
            .O(N__20695),
            .I(N__20668));
    InMux I__2105 (
            .O(N__20692),
            .I(N__20668));
    InMux I__2104 (
            .O(N__20691),
            .I(N__20665));
    InMux I__2103 (
            .O(N__20690),
            .I(N__20660));
    InMux I__2102 (
            .O(N__20689),
            .I(N__20660));
    LocalMux I__2101 (
            .O(N__20686),
            .I(N__20655));
    LocalMux I__2100 (
            .O(N__20683),
            .I(N__20655));
    LocalMux I__2099 (
            .O(N__20678),
            .I(N__20652));
    Span4Mux_v I__2098 (
            .O(N__20675),
            .I(N__20645));
    LocalMux I__2097 (
            .O(N__20668),
            .I(N__20645));
    LocalMux I__2096 (
            .O(N__20665),
            .I(N__20645));
    LocalMux I__2095 (
            .O(N__20660),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv12 I__2094 (
            .O(N__20655),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__2093 (
            .O(N__20652),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__2092 (
            .O(N__20645),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__2091 (
            .O(N__20636),
            .I(N__20633));
    LocalMux I__2090 (
            .O(N__20633),
            .I(N__20629));
    InMux I__2089 (
            .O(N__20632),
            .I(N__20626));
    Span4Mux_v I__2088 (
            .O(N__20629),
            .I(N__20623));
    LocalMux I__2087 (
            .O(N__20626),
            .I(N__20620));
    Odrv4 I__2086 (
            .O(N__20623),
            .I(\pwm_generator_inst.un3_threshold ));
    Odrv4 I__2085 (
            .O(N__20620),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__2084 (
            .O(N__20615),
            .I(N__20612));
    LocalMux I__2083 (
            .O(N__20612),
            .I(N__20609));
    Span4Mux_v I__2082 (
            .O(N__20609),
            .I(N__20606));
    Odrv4 I__2081 (
            .O(N__20606),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__2080 (
            .O(N__20603),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    CascadeMux I__2079 (
            .O(N__20600),
            .I(N__20597));
    InMux I__2078 (
            .O(N__20597),
            .I(N__20593));
    InMux I__2077 (
            .O(N__20596),
            .I(N__20590));
    LocalMux I__2076 (
            .O(N__20593),
            .I(N__20585));
    LocalMux I__2075 (
            .O(N__20590),
            .I(N__20585));
    Span4Mux_h I__2074 (
            .O(N__20585),
            .I(N__20582));
    Odrv4 I__2073 (
            .O(N__20582),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__2072 (
            .O(N__20579),
            .I(N__20575));
    InMux I__2071 (
            .O(N__20578),
            .I(N__20572));
    LocalMux I__2070 (
            .O(N__20575),
            .I(N__20569));
    LocalMux I__2069 (
            .O(N__20572),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    Odrv4 I__2068 (
            .O(N__20569),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    CascadeMux I__2067 (
            .O(N__20564),
            .I(N__20557));
    CascadeMux I__2066 (
            .O(N__20563),
            .I(N__20554));
    CascadeMux I__2065 (
            .O(N__20562),
            .I(N__20550));
    CascadeMux I__2064 (
            .O(N__20561),
            .I(N__20547));
    CascadeMux I__2063 (
            .O(N__20560),
            .I(N__20544));
    InMux I__2062 (
            .O(N__20557),
            .I(N__20533));
    InMux I__2061 (
            .O(N__20554),
            .I(N__20533));
    InMux I__2060 (
            .O(N__20553),
            .I(N__20533));
    InMux I__2059 (
            .O(N__20550),
            .I(N__20533));
    InMux I__2058 (
            .O(N__20547),
            .I(N__20533));
    InMux I__2057 (
            .O(N__20544),
            .I(N__20526));
    LocalMux I__2056 (
            .O(N__20533),
            .I(N__20523));
    InMux I__2055 (
            .O(N__20532),
            .I(N__20514));
    InMux I__2054 (
            .O(N__20531),
            .I(N__20514));
    InMux I__2053 (
            .O(N__20530),
            .I(N__20514));
    InMux I__2052 (
            .O(N__20529),
            .I(N__20514));
    LocalMux I__2051 (
            .O(N__20526),
            .I(N__20507));
    Span4Mux_h I__2050 (
            .O(N__20523),
            .I(N__20507));
    LocalMux I__2049 (
            .O(N__20514),
            .I(N__20507));
    Odrv4 I__2048 (
            .O(N__20507),
            .I(\pwm_generator_inst.N_16 ));
    InMux I__2047 (
            .O(N__20504),
            .I(N__20500));
    InMux I__2046 (
            .O(N__20503),
            .I(N__20497));
    LocalMux I__2045 (
            .O(N__20500),
            .I(N__20494));
    LocalMux I__2044 (
            .O(N__20497),
            .I(N__20491));
    Odrv4 I__2043 (
            .O(N__20494),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    Odrv4 I__2042 (
            .O(N__20491),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__2041 (
            .O(N__20486),
            .I(N__20483));
    LocalMux I__2040 (
            .O(N__20483),
            .I(N__20480));
    Span4Mux_v I__2039 (
            .O(N__20480),
            .I(N__20477));
    Odrv4 I__2038 (
            .O(N__20477),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__2037 (
            .O(N__20474),
            .I(N__20471));
    LocalMux I__2036 (
            .O(N__20471),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__2035 (
            .O(N__20468),
            .I(N__20465));
    LocalMux I__2034 (
            .O(N__20465),
            .I(N__20462));
    Span4Mux_h I__2033 (
            .O(N__20462),
            .I(N__20459));
    Odrv4 I__2032 (
            .O(N__20459),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__2031 (
            .O(N__20456),
            .I(N__20453));
    LocalMux I__2030 (
            .O(N__20453),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__2029 (
            .O(N__20450),
            .I(N__20447));
    LocalMux I__2028 (
            .O(N__20447),
            .I(N__20444));
    Span4Mux_v I__2027 (
            .O(N__20444),
            .I(N__20441));
    Odrv4 I__2026 (
            .O(N__20441),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__2025 (
            .O(N__20438),
            .I(N__20435));
    LocalMux I__2024 (
            .O(N__20435),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__2023 (
            .O(N__20432),
            .I(N__20429));
    LocalMux I__2022 (
            .O(N__20429),
            .I(N__20426));
    Span4Mux_v I__2021 (
            .O(N__20426),
            .I(N__20423));
    Odrv4 I__2020 (
            .O(N__20423),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__2019 (
            .O(N__20420),
            .I(N__20417));
    LocalMux I__2018 (
            .O(N__20417),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    CascadeMux I__2017 (
            .O(N__20414),
            .I(N__20411));
    InMux I__2016 (
            .O(N__20411),
            .I(N__20408));
    LocalMux I__2015 (
            .O(N__20408),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ));
    InMux I__2014 (
            .O(N__20405),
            .I(N__20402));
    LocalMux I__2013 (
            .O(N__20402),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ));
    InMux I__2012 (
            .O(N__20399),
            .I(N__20396));
    LocalMux I__2011 (
            .O(N__20396),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ));
    CascadeMux I__2010 (
            .O(N__20393),
            .I(N__20390));
    InMux I__2009 (
            .O(N__20390),
            .I(N__20387));
    LocalMux I__2008 (
            .O(N__20387),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ));
    InMux I__2007 (
            .O(N__20384),
            .I(N__20381));
    LocalMux I__2006 (
            .O(N__20381),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ));
    InMux I__2005 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__2004 (
            .O(N__20375),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ));
    InMux I__2003 (
            .O(N__20372),
            .I(N__20369));
    LocalMux I__2002 (
            .O(N__20369),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ));
    CascadeMux I__2001 (
            .O(N__20366),
            .I(N__20358));
    CascadeMux I__2000 (
            .O(N__20365),
            .I(N__20354));
    CascadeMux I__1999 (
            .O(N__20364),
            .I(N__20351));
    InMux I__1998 (
            .O(N__20363),
            .I(N__20346));
    InMux I__1997 (
            .O(N__20362),
            .I(N__20346));
    InMux I__1996 (
            .O(N__20361),
            .I(N__20340));
    InMux I__1995 (
            .O(N__20358),
            .I(N__20310));
    InMux I__1994 (
            .O(N__20357),
            .I(N__20310));
    InMux I__1993 (
            .O(N__20354),
            .I(N__20310));
    InMux I__1992 (
            .O(N__20351),
            .I(N__20310));
    LocalMux I__1991 (
            .O(N__20346),
            .I(N__20307));
    InMux I__1990 (
            .O(N__20345),
            .I(N__20300));
    InMux I__1989 (
            .O(N__20344),
            .I(N__20300));
    InMux I__1988 (
            .O(N__20343),
            .I(N__20300));
    LocalMux I__1987 (
            .O(N__20340),
            .I(N__20297));
    InMux I__1986 (
            .O(N__20339),
            .I(N__20286));
    InMux I__1985 (
            .O(N__20338),
            .I(N__20286));
    InMux I__1984 (
            .O(N__20337),
            .I(N__20286));
    InMux I__1983 (
            .O(N__20336),
            .I(N__20286));
    InMux I__1982 (
            .O(N__20335),
            .I(N__20286));
    InMux I__1981 (
            .O(N__20334),
            .I(N__20268));
    InMux I__1980 (
            .O(N__20333),
            .I(N__20268));
    InMux I__1979 (
            .O(N__20332),
            .I(N__20268));
    InMux I__1978 (
            .O(N__20331),
            .I(N__20268));
    InMux I__1977 (
            .O(N__20330),
            .I(N__20268));
    InMux I__1976 (
            .O(N__20329),
            .I(N__20268));
    InMux I__1975 (
            .O(N__20328),
            .I(N__20268));
    InMux I__1974 (
            .O(N__20327),
            .I(N__20268));
    InMux I__1973 (
            .O(N__20326),
            .I(N__20253));
    InMux I__1972 (
            .O(N__20325),
            .I(N__20253));
    InMux I__1971 (
            .O(N__20324),
            .I(N__20253));
    InMux I__1970 (
            .O(N__20323),
            .I(N__20253));
    InMux I__1969 (
            .O(N__20322),
            .I(N__20253));
    InMux I__1968 (
            .O(N__20321),
            .I(N__20253));
    InMux I__1967 (
            .O(N__20320),
            .I(N__20253));
    CascadeMux I__1966 (
            .O(N__20319),
            .I(N__20250));
    LocalMux I__1965 (
            .O(N__20310),
            .I(N__20247));
    Span4Mux_s1_h I__1964 (
            .O(N__20307),
            .I(N__20242));
    LocalMux I__1963 (
            .O(N__20300),
            .I(N__20242));
    Span4Mux_v I__1962 (
            .O(N__20297),
            .I(N__20237));
    LocalMux I__1961 (
            .O(N__20286),
            .I(N__20237));
    InMux I__1960 (
            .O(N__20285),
            .I(N__20234));
    LocalMux I__1959 (
            .O(N__20268),
            .I(N__20229));
    LocalMux I__1958 (
            .O(N__20253),
            .I(N__20229));
    InMux I__1957 (
            .O(N__20250),
            .I(N__20226));
    Span4Mux_h I__1956 (
            .O(N__20247),
            .I(N__20221));
    Span4Mux_v I__1955 (
            .O(N__20242),
            .I(N__20221));
    Span4Mux_v I__1954 (
            .O(N__20237),
            .I(N__20218));
    LocalMux I__1953 (
            .O(N__20234),
            .I(N__20215));
    Span4Mux_s1_h I__1952 (
            .O(N__20229),
            .I(N__20212));
    LocalMux I__1951 (
            .O(N__20226),
            .I(N__20207));
    Sp12to4 I__1950 (
            .O(N__20221),
            .I(N__20207));
    Odrv4 I__1949 (
            .O(N__20218),
            .I(N_19_1));
    Odrv12 I__1948 (
            .O(N__20215),
            .I(N_19_1));
    Odrv4 I__1947 (
            .O(N__20212),
            .I(N_19_1));
    Odrv12 I__1946 (
            .O(N__20207),
            .I(N_19_1));
    InMux I__1945 (
            .O(N__20198),
            .I(N__20195));
    LocalMux I__1944 (
            .O(N__20195),
            .I(N__20191));
    InMux I__1943 (
            .O(N__20194),
            .I(N__20188));
    Span4Mux_v I__1942 (
            .O(N__20191),
            .I(N__20185));
    LocalMux I__1941 (
            .O(N__20188),
            .I(N__20182));
    Span4Mux_v I__1940 (
            .O(N__20185),
            .I(N__20179));
    Odrv4 I__1939 (
            .O(N__20182),
            .I(\pwm_generator_inst.O_10 ));
    Odrv4 I__1938 (
            .O(N__20179),
            .I(\pwm_generator_inst.O_10 ));
    CascadeMux I__1937 (
            .O(N__20174),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__1936 (
            .O(N__20171),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__1935 (
            .O(N__20168),
            .I(N__20150));
    InMux I__1934 (
            .O(N__20167),
            .I(N__20150));
    InMux I__1933 (
            .O(N__20166),
            .I(N__20150));
    InMux I__1932 (
            .O(N__20165),
            .I(N__20150));
    InMux I__1931 (
            .O(N__20164),
            .I(N__20145));
    InMux I__1930 (
            .O(N__20163),
            .I(N__20145));
    InMux I__1929 (
            .O(N__20162),
            .I(N__20136));
    InMux I__1928 (
            .O(N__20161),
            .I(N__20136));
    InMux I__1927 (
            .O(N__20160),
            .I(N__20136));
    InMux I__1926 (
            .O(N__20159),
            .I(N__20136));
    LocalMux I__1925 (
            .O(N__20150),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__1924 (
            .O(N__20145),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__1923 (
            .O(N__20136),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__1922 (
            .O(N__20129),
            .I(N__20126));
    LocalMux I__1921 (
            .O(N__20126),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ));
    CascadeMux I__1920 (
            .O(N__20123),
            .I(N__20120));
    InMux I__1919 (
            .O(N__20120),
            .I(N__20116));
    InMux I__1918 (
            .O(N__20119),
            .I(N__20113));
    LocalMux I__1917 (
            .O(N__20116),
            .I(N__20108));
    LocalMux I__1916 (
            .O(N__20113),
            .I(N__20108));
    Span4Mux_v I__1915 (
            .O(N__20108),
            .I(N__20105));
    Odrv4 I__1914 (
            .O(N__20105),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__1913 (
            .O(N__20102),
            .I(N__20099));
    LocalMux I__1912 (
            .O(N__20099),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ));
    InMux I__1911 (
            .O(N__20096),
            .I(N__20093));
    LocalMux I__1910 (
            .O(N__20093),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__1909 (
            .O(N__20090),
            .I(N__20087));
    LocalMux I__1908 (
            .O(N__20087),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ));
    InMux I__1907 (
            .O(N__20084),
            .I(N__20081));
    LocalMux I__1906 (
            .O(N__20081),
            .I(N__20078));
    Odrv12 I__1905 (
            .O(N__20078),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__1904 (
            .O(N__20075),
            .I(N__20072));
    LocalMux I__1903 (
            .O(N__20072),
            .I(N__20069));
    Odrv12 I__1902 (
            .O(N__20069),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__1901 (
            .O(N__20066),
            .I(N__20063));
    LocalMux I__1900 (
            .O(N__20063),
            .I(N__20060));
    Odrv12 I__1899 (
            .O(N__20060),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__1898 (
            .O(N__20057),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__1897 (
            .O(N__20054),
            .I(N__20051));
    LocalMux I__1896 (
            .O(N__20051),
            .I(N__20048));
    Odrv4 I__1895 (
            .O(N__20048),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__1894 (
            .O(N__20045),
            .I(N__20042));
    LocalMux I__1893 (
            .O(N__20042),
            .I(N_86_i_i));
    InMux I__1892 (
            .O(N__20039),
            .I(bfn_1_23_0_));
    InMux I__1891 (
            .O(N__20036),
            .I(N__20033));
    LocalMux I__1890 (
            .O(N__20033),
            .I(N__20030));
    Span4Mux_v I__1889 (
            .O(N__20030),
            .I(N__20027));
    Odrv4 I__1888 (
            .O(N__20027),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__1887 (
            .O(N__20024),
            .I(N__20021));
    LocalMux I__1886 (
            .O(N__20021),
            .I(N__20018));
    Odrv12 I__1885 (
            .O(N__20018),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__1884 (
            .O(N__20015),
            .I(N__20012));
    LocalMux I__1883 (
            .O(N__20012),
            .I(N__20009));
    Odrv12 I__1882 (
            .O(N__20009),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__1881 (
            .O(N__20006),
            .I(N__20003));
    LocalMux I__1880 (
            .O(N__20003),
            .I(N__20000));
    Odrv12 I__1879 (
            .O(N__20000),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__1878 (
            .O(N__19997),
            .I(N__19994));
    LocalMux I__1877 (
            .O(N__19994),
            .I(N__19991));
    Odrv12 I__1876 (
            .O(N__19991),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__1875 (
            .O(N__19988),
            .I(N__19985));
    LocalMux I__1874 (
            .O(N__19985),
            .I(N__19982));
    Odrv4 I__1873 (
            .O(N__19982),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__1872 (
            .O(N__19979),
            .I(N__19976));
    LocalMux I__1871 (
            .O(N__19976),
            .I(N__19973));
    Odrv4 I__1870 (
            .O(N__19973),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__1869 (
            .O(N__19970),
            .I(N__19967));
    LocalMux I__1868 (
            .O(N__19967),
            .I(N__19964));
    Odrv12 I__1867 (
            .O(N__19964),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__1866 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__1865 (
            .O(N__19958),
            .I(N__19955));
    Odrv4 I__1864 (
            .O(N__19955),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1863 (
            .O(N__19952),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__1862 (
            .O(N__19949),
            .I(N__19946));
    LocalMux I__1861 (
            .O(N__19946),
            .I(N__19943));
    Odrv4 I__1860 (
            .O(N__19943),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1859 (
            .O(N__19940),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__1858 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__1857 (
            .O(N__19934),
            .I(N__19931));
    Odrv4 I__1856 (
            .O(N__19931),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1855 (
            .O(N__19928),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__1854 (
            .O(N__19925),
            .I(N__19922));
    LocalMux I__1853 (
            .O(N__19922),
            .I(N__19919));
    Span4Mux_v I__1852 (
            .O(N__19919),
            .I(N__19916));
    Odrv4 I__1851 (
            .O(N__19916),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__1850 (
            .O(N__19913),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    CascadeMux I__1849 (
            .O(N__19910),
            .I(N__19907));
    InMux I__1848 (
            .O(N__19907),
            .I(N__19904));
    LocalMux I__1847 (
            .O(N__19904),
            .I(N__19901));
    Odrv12 I__1846 (
            .O(N__19901),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__1845 (
            .O(N__19898),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__1844 (
            .O(N__19895),
            .I(N__19892));
    LocalMux I__1843 (
            .O(N__19892),
            .I(N__19889));
    Odrv4 I__1842 (
            .O(N__19889),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__1841 (
            .O(N__19886),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    CascadeMux I__1840 (
            .O(N__19883),
            .I(N__19880));
    InMux I__1839 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__1838 (
            .O(N__19877),
            .I(N__19874));
    Odrv4 I__1837 (
            .O(N__19874),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__1836 (
            .O(N__19871),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__1835 (
            .O(N__19868),
            .I(N__19865));
    LocalMux I__1834 (
            .O(N__19865),
            .I(N__19862));
    Span4Mux_v I__1833 (
            .O(N__19862),
            .I(N__19859));
    Odrv4 I__1832 (
            .O(N__19859),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__1831 (
            .O(N__19856),
            .I(N__19853));
    LocalMux I__1830 (
            .O(N__19853),
            .I(N__19850));
    Span4Mux_v I__1829 (
            .O(N__19850),
            .I(N__19847));
    Odrv4 I__1828 (
            .O(N__19847),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    InMux I__1827 (
            .O(N__19844),
            .I(N__19841));
    LocalMux I__1826 (
            .O(N__19841),
            .I(N__19838));
    Span4Mux_v I__1825 (
            .O(N__19838),
            .I(N__19835));
    Span4Mux_v I__1824 (
            .O(N__19835),
            .I(N__19832));
    Span4Mux_v I__1823 (
            .O(N__19832),
            .I(N__19829));
    Odrv4 I__1822 (
            .O(N__19829),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__1821 (
            .O(N__19826),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    InMux I__1820 (
            .O(N__19823),
            .I(N__19820));
    LocalMux I__1819 (
            .O(N__19820),
            .I(N__19817));
    Span4Mux_v I__1818 (
            .O(N__19817),
            .I(N__19813));
    InMux I__1817 (
            .O(N__19816),
            .I(N__19810));
    Span4Mux_v I__1816 (
            .O(N__19813),
            .I(N__19802));
    LocalMux I__1815 (
            .O(N__19810),
            .I(N__19802));
    CascadeMux I__1814 (
            .O(N__19809),
            .I(N__19798));
    CascadeMux I__1813 (
            .O(N__19808),
            .I(N__19794));
    CascadeMux I__1812 (
            .O(N__19807),
            .I(N__19790));
    Span4Mux_v I__1811 (
            .O(N__19802),
            .I(N__19787));
    InMux I__1810 (
            .O(N__19801),
            .I(N__19774));
    InMux I__1809 (
            .O(N__19798),
            .I(N__19774));
    InMux I__1808 (
            .O(N__19797),
            .I(N__19774));
    InMux I__1807 (
            .O(N__19794),
            .I(N__19774));
    InMux I__1806 (
            .O(N__19793),
            .I(N__19774));
    InMux I__1805 (
            .O(N__19790),
            .I(N__19774));
    Span4Mux_v I__1804 (
            .O(N__19787),
            .I(N__19769));
    LocalMux I__1803 (
            .O(N__19774),
            .I(N__19769));
    Span4Mux_v I__1802 (
            .O(N__19769),
            .I(N__19766));
    Odrv4 I__1801 (
            .O(N__19766),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    CascadeMux I__1800 (
            .O(N__19763),
            .I(N__19760));
    InMux I__1799 (
            .O(N__19760),
            .I(N__19757));
    LocalMux I__1798 (
            .O(N__19757),
            .I(N__19754));
    Span12Mux_v I__1797 (
            .O(N__19754),
            .I(N__19751));
    Odrv12 I__1796 (
            .O(N__19751),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__1795 (
            .O(N__19748),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__1794 (
            .O(N__19745),
            .I(N__19742));
    LocalMux I__1793 (
            .O(N__19742),
            .I(N__19739));
    Odrv12 I__1792 (
            .O(N__19739),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__1791 (
            .O(N__19736),
            .I(bfn_1_21_0_));
    CascadeMux I__1790 (
            .O(N__19733),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_ ));
    InMux I__1789 (
            .O(N__19730),
            .I(N__19727));
    LocalMux I__1788 (
            .O(N__19727),
            .I(N__19724));
    Span4Mux_v I__1787 (
            .O(N__19724),
            .I(N__19721));
    Odrv4 I__1786 (
            .O(N__19721),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    InMux I__1785 (
            .O(N__19718),
            .I(N__19715));
    LocalMux I__1784 (
            .O(N__19715),
            .I(N__19712));
    Odrv12 I__1783 (
            .O(N__19712),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__1782 (
            .O(N__19709),
            .I(N__19706));
    LocalMux I__1781 (
            .O(N__19706),
            .I(N__19703));
    Odrv12 I__1780 (
            .O(N__19703),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__1779 (
            .O(N__19700),
            .I(N__19697));
    LocalMux I__1778 (
            .O(N__19697),
            .I(N__19694));
    Span4Mux_s2_h I__1777 (
            .O(N__19694),
            .I(N__19691));
    Odrv4 I__1776 (
            .O(N__19691),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__1775 (
            .O(N__19688),
            .I(N__19685));
    LocalMux I__1774 (
            .O(N__19685),
            .I(N__19682));
    Odrv4 I__1773 (
            .O(N__19682),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__1772 (
            .O(N__19679),
            .I(N__19676));
    LocalMux I__1771 (
            .O(N__19676),
            .I(N__19673));
    Odrv12 I__1770 (
            .O(N__19673),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    InMux I__1769 (
            .O(N__19670),
            .I(N__19667));
    LocalMux I__1768 (
            .O(N__19667),
            .I(N__19664));
    Span4Mux_v I__1767 (
            .O(N__19664),
            .I(N__19661));
    Span4Mux_v I__1766 (
            .O(N__19661),
            .I(N__19658));
    Span4Mux_v I__1765 (
            .O(N__19658),
            .I(N__19655));
    Odrv4 I__1764 (
            .O(N__19655),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    CascadeMux I__1763 (
            .O(N__19652),
            .I(N__19649));
    InMux I__1762 (
            .O(N__19649),
            .I(N__19646));
    LocalMux I__1761 (
            .O(N__19646),
            .I(N__19643));
    Span4Mux_v I__1760 (
            .O(N__19643),
            .I(N__19640));
    Odrv4 I__1759 (
            .O(N__19640),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    InMux I__1758 (
            .O(N__19637),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__1757 (
            .O(N__19634),
            .I(N__19631));
    LocalMux I__1756 (
            .O(N__19631),
            .I(N__19628));
    Span4Mux_v I__1755 (
            .O(N__19628),
            .I(N__19625));
    Span4Mux_v I__1754 (
            .O(N__19625),
            .I(N__19622));
    Span4Mux_v I__1753 (
            .O(N__19622),
            .I(N__19619));
    Odrv4 I__1752 (
            .O(N__19619),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    CascadeMux I__1751 (
            .O(N__19616),
            .I(N__19613));
    InMux I__1750 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__1749 (
            .O(N__19610),
            .I(N__19607));
    Span4Mux_v I__1748 (
            .O(N__19607),
            .I(N__19604));
    Odrv4 I__1747 (
            .O(N__19604),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    InMux I__1746 (
            .O(N__19601),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__1745 (
            .O(N__19598),
            .I(N__19595));
    LocalMux I__1744 (
            .O(N__19595),
            .I(N__19592));
    Span4Mux_v I__1743 (
            .O(N__19592),
            .I(N__19589));
    Span4Mux_v I__1742 (
            .O(N__19589),
            .I(N__19586));
    Span4Mux_v I__1741 (
            .O(N__19586),
            .I(N__19583));
    Odrv4 I__1740 (
            .O(N__19583),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    CascadeMux I__1739 (
            .O(N__19580),
            .I(N__19577));
    InMux I__1738 (
            .O(N__19577),
            .I(N__19574));
    LocalMux I__1737 (
            .O(N__19574),
            .I(N__19571));
    Span4Mux_v I__1736 (
            .O(N__19571),
            .I(N__19568));
    Odrv4 I__1735 (
            .O(N__19568),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    InMux I__1734 (
            .O(N__19565),
            .I(bfn_1_20_0_));
    InMux I__1733 (
            .O(N__19562),
            .I(N__19559));
    LocalMux I__1732 (
            .O(N__19559),
            .I(N__19556));
    Span4Mux_v I__1731 (
            .O(N__19556),
            .I(N__19553));
    Span4Mux_v I__1730 (
            .O(N__19553),
            .I(N__19550));
    Span4Mux_v I__1729 (
            .O(N__19550),
            .I(N__19547));
    Odrv4 I__1728 (
            .O(N__19547),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    CascadeMux I__1727 (
            .O(N__19544),
            .I(N__19541));
    InMux I__1726 (
            .O(N__19541),
            .I(N__19538));
    LocalMux I__1725 (
            .O(N__19538),
            .I(N__19535));
    Span4Mux_v I__1724 (
            .O(N__19535),
            .I(N__19532));
    Odrv4 I__1723 (
            .O(N__19532),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    InMux I__1722 (
            .O(N__19529),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    InMux I__1721 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__1720 (
            .O(N__19523),
            .I(N__19520));
    Span12Mux_h I__1719 (
            .O(N__19520),
            .I(N__19517));
    Span12Mux_v I__1718 (
            .O(N__19517),
            .I(N__19514));
    Odrv12 I__1717 (
            .O(N__19514),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__1716 (
            .O(N__19511),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    CascadeMux I__1715 (
            .O(N__19508),
            .I(N__19505));
    InMux I__1714 (
            .O(N__19505),
            .I(N__19502));
    LocalMux I__1713 (
            .O(N__19502),
            .I(N__19499));
    Span4Mux_h I__1712 (
            .O(N__19499),
            .I(N__19496));
    Span4Mux_v I__1711 (
            .O(N__19496),
            .I(N__19493));
    Sp12to4 I__1710 (
            .O(N__19493),
            .I(N__19490));
    Odrv12 I__1709 (
            .O(N__19490),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__1708 (
            .O(N__19487),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    InMux I__1707 (
            .O(N__19484),
            .I(N__19481));
    LocalMux I__1706 (
            .O(N__19481),
            .I(N__19478));
    Span4Mux_v I__1705 (
            .O(N__19478),
            .I(N__19475));
    Span4Mux_v I__1704 (
            .O(N__19475),
            .I(N__19472));
    Span4Mux_v I__1703 (
            .O(N__19472),
            .I(N__19469));
    Odrv4 I__1702 (
            .O(N__19469),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__1701 (
            .O(N__19466),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    CascadeMux I__1700 (
            .O(N__19463),
            .I(N__19460));
    InMux I__1699 (
            .O(N__19460),
            .I(N__19457));
    LocalMux I__1698 (
            .O(N__19457),
            .I(N__19454));
    Span4Mux_h I__1697 (
            .O(N__19454),
            .I(N__19451));
    Sp12to4 I__1696 (
            .O(N__19451),
            .I(N__19448));
    Span12Mux_v I__1695 (
            .O(N__19448),
            .I(N__19445));
    Odrv12 I__1694 (
            .O(N__19445),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__1693 (
            .O(N__19442),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    InMux I__1692 (
            .O(N__19439),
            .I(N__19436));
    LocalMux I__1691 (
            .O(N__19436),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    InMux I__1690 (
            .O(N__19433),
            .I(N__19430));
    LocalMux I__1689 (
            .O(N__19430),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__1688 (
            .O(N__19427),
            .I(N__19424));
    LocalMux I__1687 (
            .O(N__19424),
            .I(N__19421));
    Span4Mux_v I__1686 (
            .O(N__19421),
            .I(N__19418));
    Span4Mux_v I__1685 (
            .O(N__19418),
            .I(N__19415));
    Span4Mux_v I__1684 (
            .O(N__19415),
            .I(N__19412));
    Odrv4 I__1683 (
            .O(N__19412),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__1682 (
            .O(N__19409),
            .I(N__19406));
    InMux I__1681 (
            .O(N__19406),
            .I(N__19403));
    LocalMux I__1680 (
            .O(N__19403),
            .I(N__19400));
    Span4Mux_v I__1679 (
            .O(N__19400),
            .I(N__19397));
    Odrv4 I__1678 (
            .O(N__19397),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__1677 (
            .O(N__19394),
            .I(N__19391));
    LocalMux I__1676 (
            .O(N__19391),
            .I(N__19388));
    Span4Mux_v I__1675 (
            .O(N__19388),
            .I(N__19385));
    Span4Mux_v I__1674 (
            .O(N__19385),
            .I(N__19382));
    Span4Mux_v I__1673 (
            .O(N__19382),
            .I(N__19379));
    Odrv4 I__1672 (
            .O(N__19379),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__1671 (
            .O(N__19376),
            .I(N__19373));
    InMux I__1670 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__1669 (
            .O(N__19370),
            .I(N__19367));
    Span4Mux_v I__1668 (
            .O(N__19367),
            .I(N__19364));
    Odrv4 I__1667 (
            .O(N__19364),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    InMux I__1666 (
            .O(N__19361),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__1665 (
            .O(N__19358),
            .I(N__19355));
    LocalMux I__1664 (
            .O(N__19355),
            .I(N__19352));
    Span12Mux_h I__1663 (
            .O(N__19352),
            .I(N__19349));
    Span12Mux_v I__1662 (
            .O(N__19349),
            .I(N__19346));
    Odrv12 I__1661 (
            .O(N__19346),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__1660 (
            .O(N__19343),
            .I(N__19340));
    InMux I__1659 (
            .O(N__19340),
            .I(N__19337));
    LocalMux I__1658 (
            .O(N__19337),
            .I(N__19334));
    Span4Mux_v I__1657 (
            .O(N__19334),
            .I(N__19331));
    Odrv4 I__1656 (
            .O(N__19331),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__1655 (
            .O(N__19328),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__1654 (
            .O(N__19325),
            .I(N__19322));
    LocalMux I__1653 (
            .O(N__19322),
            .I(N__19319));
    Span4Mux_v I__1652 (
            .O(N__19319),
            .I(N__19316));
    Span4Mux_v I__1651 (
            .O(N__19316),
            .I(N__19313));
    Span4Mux_v I__1650 (
            .O(N__19313),
            .I(N__19310));
    Odrv4 I__1649 (
            .O(N__19310),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__1648 (
            .O(N__19307),
            .I(N__19304));
    InMux I__1647 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__1646 (
            .O(N__19301),
            .I(N__19298));
    Span4Mux_v I__1645 (
            .O(N__19298),
            .I(N__19295));
    Odrv4 I__1644 (
            .O(N__19295),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    InMux I__1643 (
            .O(N__19292),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__1642 (
            .O(N__19289),
            .I(N__19286));
    LocalMux I__1641 (
            .O(N__19286),
            .I(N__19283));
    Span4Mux_v I__1640 (
            .O(N__19283),
            .I(N__19280));
    Span4Mux_v I__1639 (
            .O(N__19280),
            .I(N__19277));
    Span4Mux_v I__1638 (
            .O(N__19277),
            .I(N__19274));
    Odrv4 I__1637 (
            .O(N__19274),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__1636 (
            .O(N__19271),
            .I(N__19268));
    InMux I__1635 (
            .O(N__19268),
            .I(N__19265));
    LocalMux I__1634 (
            .O(N__19265),
            .I(N__19262));
    Span4Mux_v I__1633 (
            .O(N__19262),
            .I(N__19259));
    Span4Mux_v I__1632 (
            .O(N__19259),
            .I(N__19256));
    Odrv4 I__1631 (
            .O(N__19256),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__1630 (
            .O(N__19253),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__1629 (
            .O(N__19250),
            .I(N__19247));
    LocalMux I__1628 (
            .O(N__19247),
            .I(N__19244));
    Span4Mux_v I__1627 (
            .O(N__19244),
            .I(N__19241));
    Span4Mux_v I__1626 (
            .O(N__19241),
            .I(N__19238));
    Span4Mux_v I__1625 (
            .O(N__19238),
            .I(N__19235));
    Odrv4 I__1624 (
            .O(N__19235),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__1623 (
            .O(N__19232),
            .I(N__19229));
    InMux I__1622 (
            .O(N__19229),
            .I(N__19226));
    LocalMux I__1621 (
            .O(N__19226),
            .I(N__19223));
    Span4Mux_h I__1620 (
            .O(N__19223),
            .I(N__19220));
    Span4Mux_v I__1619 (
            .O(N__19220),
            .I(N__19217));
    Odrv4 I__1618 (
            .O(N__19217),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__1617 (
            .O(N__19214),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__1616 (
            .O(N__19211),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    InMux I__1615 (
            .O(N__19208),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__1614 (
            .O(N__19205),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__1613 (
            .O(N__19202),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__1612 (
            .O(N__19199),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__1611 (
            .O(N__19196),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__1610 (
            .O(N__19193),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    InMux I__1609 (
            .O(N__19190),
            .I(bfn_1_18_0_));
    InMux I__1608 (
            .O(N__19187),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    InMux I__1607 (
            .O(N__19184),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__1606 (
            .O(N__19181),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__1605 (
            .O(N__19178),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__1604 (
            .O(N__19175),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__1603 (
            .O(N__19172),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__1602 (
            .O(N__19169),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__1601 (
            .O(N__19166),
            .I(bfn_1_16_0_));
    InMux I__1600 (
            .O(N__19163),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__1599 (
            .O(N__19160),
            .I(N__19157));
    LocalMux I__1598 (
            .O(N__19157),
            .I(N__19154));
    Span4Mux_v I__1597 (
            .O(N__19154),
            .I(N__19150));
    InMux I__1596 (
            .O(N__19153),
            .I(N__19147));
    Odrv4 I__1595 (
            .O(N__19150),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    LocalMux I__1594 (
            .O(N__19147),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    InMux I__1593 (
            .O(N__19142),
            .I(N__19139));
    LocalMux I__1592 (
            .O(N__19139),
            .I(N__19136));
    Span4Mux_v I__1591 (
            .O(N__19136),
            .I(N__19133));
    Odrv4 I__1590 (
            .O(N__19133),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__1589 (
            .O(N__19130),
            .I(bfn_1_15_0_));
    InMux I__1588 (
            .O(N__19127),
            .I(\pwm_generator_inst.counter_cry_0 ));
    IoInMux I__1587 (
            .O(N__19124),
            .I(N__19121));
    LocalMux I__1586 (
            .O(N__19121),
            .I(N__19118));
    Span4Mux_s3_v I__1585 (
            .O(N__19118),
            .I(N__19115));
    Span4Mux_h I__1584 (
            .O(N__19115),
            .I(N__19112));
    Sp12to4 I__1583 (
            .O(N__19112),
            .I(N__19109));
    Span12Mux_v I__1582 (
            .O(N__19109),
            .I(N__19106));
    Span12Mux_v I__1581 (
            .O(N__19106),
            .I(N__19103));
    Odrv12 I__1580 (
            .O(N__19103),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1579 (
            .O(N__19100),
            .I(N__19097));
    LocalMux I__1578 (
            .O(N__19097),
            .I(N__19094));
    IoSpan4Mux I__1577 (
            .O(N__19094),
            .I(N__19091));
    IoSpan4Mux I__1576 (
            .O(N__19091),
            .I(N__19088));
    Odrv4 I__1575 (
            .O(N__19088),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_15_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_5_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_15_6_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_5_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_19_0_));
    defparam IN_MUX_bfv_5_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_5_20_0_));
    defparam IN_MUX_bfv_5_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_21_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_5_21_0_));
    defparam IN_MUX_bfv_5_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_22_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_5_22_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_2_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_21_0_));
    defparam IN_MUX_bfv_2_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_22_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_2_22_0_));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_14_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_4_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_18_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_7_0_));
    defparam IN_MUX_bfv_18_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_8_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_15 ),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_23 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_18_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_22_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_18_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_23_0_));
    defparam IN_MUX_bfv_18_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_18_24_0_));
    defparam IN_MUX_bfv_18_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_25_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_18_25_0_));
    defparam IN_MUX_bfv_18_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_26_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_18_26_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_11_22_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19124),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19100),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__35834),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_161_i_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__26210),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__36881),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__44747),
            .CLKHFEN(N__44786),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__44785),
            .RGB2PWM(N__20045),
            .RGB1(rgb_g),
            .CURREN(N__44831),
            .RGB2(rgb_b),
            .RGB1PWM(N__21068),
            .RGB0PWM(N__49271),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_6_3  (
            .in0(N__19823),
            .in1(N__19153),
            .in2(_gnd_net_),
            .in3(N__20285),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25250),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50049),
            .ce(),
            .sr(N__49207));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_1  (
            .in0(N__19160),
            .in1(N__19816),
            .in2(N__20319),
            .in3(N__19142),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_1_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_1_15_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_1_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_1_15_0  (
            .in0(N__20165),
            .in1(N__21238),
            .in2(_gnd_net_),
            .in3(N__19130),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__50020),
            .ce(),
            .sr(N__49227));
    defparam \pwm_generator_inst.counter_1_LC_1_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_1_15_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_1_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_1_15_1  (
            .in0(N__20159),
            .in1(N__21196),
            .in2(_gnd_net_),
            .in3(N__19127),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__50020),
            .ce(),
            .sr(N__49227));
    defparam \pwm_generator_inst.counter_2_LC_1_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_1_15_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_1_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_1_15_2  (
            .in0(N__20166),
            .in1(N__21520),
            .in2(_gnd_net_),
            .in3(N__19184),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__50020),
            .ce(),
            .sr(N__49227));
    defparam \pwm_generator_inst.counter_3_LC_1_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_1_15_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_1_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_1_15_3  (
            .in0(N__20160),
            .in1(N__21493),
            .in2(_gnd_net_),
            .in3(N__19181),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__50020),
            .ce(),
            .sr(N__49227));
    defparam \pwm_generator_inst.counter_4_LC_1_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_1_15_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_1_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_1_15_4  (
            .in0(N__20167),
            .in1(N__21448),
            .in2(_gnd_net_),
            .in3(N__19178),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__50020),
            .ce(),
            .sr(N__49227));
    defparam \pwm_generator_inst.counter_5_LC_1_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_1_15_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_1_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_1_15_5  (
            .in0(N__20161),
            .in1(N__21396),
            .in2(_gnd_net_),
            .in3(N__19175),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__50020),
            .ce(),
            .sr(N__49227));
    defparam \pwm_generator_inst.counter_6_LC_1_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_1_15_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_1_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_1_15_6  (
            .in0(N__20168),
            .in1(N__21357),
            .in2(_gnd_net_),
            .in3(N__19172),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__50020),
            .ce(),
            .sr(N__49227));
    defparam \pwm_generator_inst.counter_7_LC_1_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_1_15_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_1_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_1_15_7  (
            .in0(N__20162),
            .in1(N__21319),
            .in2(_gnd_net_),
            .in3(N__19169),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__50020),
            .ce(),
            .sr(N__49227));
    defparam \pwm_generator_inst.counter_8_LC_1_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_1_16_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_1_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_1_16_0  (
            .in0(N__20164),
            .in1(N__21280),
            .in2(_gnd_net_),
            .in3(N__19166),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__50010),
            .ce(),
            .sr(N__49233));
    defparam \pwm_generator_inst.counter_9_LC_1_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_1_16_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_1_16_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_1_16_1  (
            .in0(N__21649),
            .in1(N__20163),
            .in2(_gnd_net_),
            .in3(N__19163),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50010),
            .ce(),
            .sr(N__49233));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_1_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_1_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__19730),
            .in2(N__20713),
            .in3(N__20707),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_1_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_1_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__20615),
            .in2(_gnd_net_),
            .in3(N__19211),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_1_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_1_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__19439),
            .in2(_gnd_net_),
            .in3(N__19208),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_1_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_1_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__19433),
            .in2(_gnd_net_),
            .in3(N__19205),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_1_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_1_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__19718),
            .in2(_gnd_net_),
            .in3(N__19202),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_1_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_1_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__19709),
            .in2(_gnd_net_),
            .in3(N__19199),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_1_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_1_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__19700),
            .in2(_gnd_net_),
            .in3(N__19196),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_1_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_1_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__19679),
            .in2(_gnd_net_),
            .in3(N__19193),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_1_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_1_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__19688),
            .in2(_gnd_net_),
            .in3(N__19190),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_1_18_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_1_18_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_1_18_1  (
            .in0(N__20867),
            .in1(N__19856),
            .in2(N__20714),
            .in3(N__19187),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_1_18_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_1_18_5 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_1_18_5  (
            .in0(N__21035),
            .in1(N__21054),
            .in2(N__20600),
            .in3(N__20702),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_1_18_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_1_18_6 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_1_18_6  (
            .in0(N__20703),
            .in1(N__21020),
            .in2(N__20123),
            .in3(N__20996),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_19_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__19427),
            .in2(N__19409),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_1_19_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_1_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__19394),
            .in2(N__19376),
            .in3(N__19361),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_1_19_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_1_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__19358),
            .in2(N__19343),
            .in3(N__19328),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_1_19_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_1_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(N__19325),
            .in2(N__19307),
            .in3(N__19292),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_1_19_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_1_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(N__19289),
            .in2(N__19271),
            .in3(N__19253),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_1_19_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_1_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__19250),
            .in2(N__19232),
            .in3(N__19214),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_1_19_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_1_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(N__19670),
            .in2(N__19652),
            .in3(N__19637),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_1_19_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_1_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__19634),
            .in2(N__19616),
            .in3(N__19601),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_1_20_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_1_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(N__19598),
            .in2(N__19580),
            .in3(N__19565),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_1_20_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_1_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__19562),
            .in2(N__19544),
            .in3(N__19529),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_1_20_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_1_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(N__19526),
            .in2(N__19807),
            .in3(N__19511),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_1_20_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_1_20_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_1_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_1_20_3  (
            .in0(_gnd_net_),
            .in1(N__19793),
            .in2(N__19508),
            .in3(N__19487),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_1_20_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_1_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(N__19484),
            .in2(N__19808),
            .in3(N__19466),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_1_20_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_1_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_1_20_5  (
            .in0(_gnd_net_),
            .in1(N__19797),
            .in2(N__19463),
            .in3(N__19442),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_1_20_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_1_20_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_1_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_1_20_6  (
            .in0(_gnd_net_),
            .in1(N__19844),
            .in2(N__19809),
            .in3(N__19826),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_1_20_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_1_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_1_20_7  (
            .in0(_gnd_net_),
            .in1(N__19801),
            .in2(N__19763),
            .in3(N__19748),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_1_21_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_1_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_1_21_0  (
            .in0(N__19745),
            .in1(N__20054),
            .in2(_gnd_net_),
            .in3(N__19736),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_1_21_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_1_21_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_1_21_1 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_1_21_1  (
            .in0(N__20723),
            .in1(N__20194),
            .in2(N__19733),
            .in3(N__20747),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_1_21_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_1_21_2 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_1_21_2  (
            .in0(N__20981),
            .in1(N__20954),
            .in2(N__20708),
            .in3(N__20504),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_1_21_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_1_21_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_1_21_3 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_1_21_3  (
            .in0(N__20578),
            .in1(N__20921),
            .in2(N__20945),
            .in3(N__20695),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_1_21_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_1_21_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_1_21_4 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_1_21_4  (
            .in0(N__20912),
            .in1(N__21164),
            .in2(N__20709),
            .in3(N__21176),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_1_21_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_1_21_5 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_1_21_5  (
            .in0(N__20690),
            .in1(N__21128),
            .in2(N__21146),
            .in3(N__20882),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_1_21_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_1_21_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_1_21_6 .LUT_INIT=16'b1011011110000100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_1_21_6  (
            .in0(N__21086),
            .in1(N__20689),
            .in2(N__20900),
            .in3(N__21098),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_22_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(N__20632),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_22_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_22_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(N__19961),
            .in2(_gnd_net_),
            .in3(N__19952),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_22_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_22_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_22_2  (
            .in0(_gnd_net_),
            .in1(N__19949),
            .in2(_gnd_net_),
            .in3(N__19940),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_22_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(N__19937),
            .in2(_gnd_net_),
            .in3(N__19928),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_22_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(N__19925),
            .in2(_gnd_net_),
            .in3(N__19913),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_22_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_22_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(N__44716),
            .in2(N__19910),
            .in3(N__19898),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_22_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_22_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(N__19895),
            .in2(N__44746),
            .in3(N__19886),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_22_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_22_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(N__44720),
            .in2(N__19883),
            .in3(N__19871),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(N__19868),
            .in2(_gnd_net_),
            .in3(N__20039),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_23_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(N__20036),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_23_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(N__20024),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_23_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_23_3  (
            .in0(_gnd_net_),
            .in1(N__20015),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_23_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(N__20006),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_23_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_23_5  (
            .in0(_gnd_net_),
            .in1(N__19997),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(N__19988),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_23_7  (
            .in0(_gnd_net_),
            .in1(N__19979),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_24_0  (
            .in0(_gnd_net_),
            .in1(N__19970),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_24_1  (
            .in0(_gnd_net_),
            .in1(N__20084),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_24_2  (
            .in0(_gnd_net_),
            .in1(N__20075),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_24_3  (
            .in0(_gnd_net_),
            .in1(N__20066),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_24_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20057),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_25_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_25_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_25_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.N_86_i_i_LC_1_30_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_86_i_i_LC_1_30_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_86_i_i_LC_1_30_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \phase_controller_inst1.N_86_i_i_LC_1_30_3  (
            .in0(N__30008),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49270),
            .lcout(N_86_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_0 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_0  (
            .in0(N__25508),
            .in1(N__23468),
            .in2(N__22316),
            .in3(N__23276),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50032),
            .ce(),
            .sr(N__49211));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_6 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_6  (
            .in0(N__25509),
            .in1(N__23469),
            .in2(N__21938),
            .in3(N__23277),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50032),
            .ce(),
            .sr(N__49211));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_14_0 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_2_14_0  (
            .in0(N__25510),
            .in1(N__23467),
            .in2(N__22160),
            .in3(N__23269),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50021),
            .ce(),
            .sr(N__49216));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_2_15_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_2_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__21516),
            .in2(_gnd_net_),
            .in3(N__21234),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_2_15_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_2_15_5 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_2_15_5  (
            .in0(N__21447),
            .in1(N__21489),
            .in2(N__20174),
            .in3(N__21195),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_2_15_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_2_15_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_2_15_6  (
            .in0(N__20096),
            .in1(N__21358),
            .in2(N__20171),
            .in3(N__21397),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_15_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_15_7  (
            .in0(N__24453),
            .in1(N__24725),
            .in2(N__24571),
            .in3(N__24678),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_2_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_2_16_1 .LUT_INIT=16'b1101110111001111;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_2_16_1  (
            .in0(N__21592),
            .in1(N__20129),
            .in2(N__20563),
            .in3(N__20338),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_16_2  (
            .in0(N__21015),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20119),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_2_16_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_2_16_3 .LUT_INIT=16'b1101110111001111;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_2_16_3  (
            .in0(N__21593),
            .in1(N__20102),
            .in2(N__20564),
            .in3(N__20339),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_2_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_2_16_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_2_16_4  (
            .in0(N__21645),
            .in1(N__21276),
            .in2(_gnd_net_),
            .in3(N__21318),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_2_16_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_2_16_5 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_2_16_5  (
            .in0(N__21590),
            .in1(N__20090),
            .in2(N__20562),
            .in3(N__20337),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_2_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_2_16_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_2_16_6  (
            .in0(N__20336),
            .in1(N__21591),
            .in2(N__20414),
            .in3(N__20553),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_2_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_2_16_7 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_2_16_7  (
            .in0(N__21589),
            .in1(N__20405),
            .in2(N__20561),
            .in3(N__20335),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_2_17_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_2_17_1 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_2_17_1  (
            .in0(N__20529),
            .in1(N__20399),
            .in2(N__20364),
            .in3(N__21585),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_2_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_2_17_2 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_2_17_2  (
            .in0(N__21587),
            .in1(N__20531),
            .in2(N__20393),
            .in3(N__20357),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_2_17_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_2_17_3 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_2_17_3  (
            .in0(N__20532),
            .in1(N__21588),
            .in2(N__20366),
            .in3(N__20384),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_2_17_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_2_17_7 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_2_17_7  (
            .in0(N__20530),
            .in1(N__20378),
            .in2(N__20365),
            .in3(N__21586),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_2_18_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_2_18_0 .LUT_INIT=16'b1101110111001111;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_2_18_0  (
            .in0(N__21584),
            .in1(N__20372),
            .in2(N__20560),
            .in3(N__20361),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__24564),
            .in2(_gnd_net_),
            .in3(N__24726),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_18_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_18_2  (
            .in0(N__24104),
            .in1(N__23847),
            .in2(_gnd_net_),
            .in3(N__23931),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_18_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_18_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__20198),
            .in2(_gnd_net_),
            .in3(N__20745),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_18_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_18_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__20596),
            .in2(_gnd_net_),
            .in3(N__21055),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_20_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_20_1  (
            .in0(N__20943),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20579),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_20_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_20_2 .LUT_INIT=16'b1100111111001101;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_2_20_2  (
            .in0(N__21744),
            .in1(N__21875),
            .in2(N__21797),
            .in3(N__21107),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_20_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_2_20_3  (
            .in0(N__20976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20503),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_21_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_21_0  (
            .in0(_gnd_net_),
            .in1(N__20474),
            .in2(_gnd_net_),
            .in3(N__20486),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_2_21_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_21_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_21_1  (
            .in0(_gnd_net_),
            .in1(N__20456),
            .in2(_gnd_net_),
            .in3(N__20468),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_21_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_21_2  (
            .in0(_gnd_net_),
            .in1(N__20438),
            .in2(_gnd_net_),
            .in3(N__20450),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_21_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_21_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_21_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_21_3  (
            .in0(N__20432),
            .in1(N__20420),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_21_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_21_4  (
            .in0(_gnd_net_),
            .in1(N__20843),
            .in2(_gnd_net_),
            .in3(N__20855),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_21_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_21_5  (
            .in0(_gnd_net_),
            .in1(N__20825),
            .in2(_gnd_net_),
            .in3(N__20837),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_21_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_21_6  (
            .in0(_gnd_net_),
            .in1(N__20807),
            .in2(_gnd_net_),
            .in3(N__20819),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_21_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_21_7  (
            .in0(_gnd_net_),
            .in1(N__20789),
            .in2(_gnd_net_),
            .in3(N__20801),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_22_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_22_0  (
            .in0(_gnd_net_),
            .in1(N__20771),
            .in2(_gnd_net_),
            .in3(N__20783),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_2_22_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_22_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_22_1  (
            .in0(_gnd_net_),
            .in1(N__20753),
            .in2(_gnd_net_),
            .in3(N__20765),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_22_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_22_2  (
            .in0(_gnd_net_),
            .in1(N__20746),
            .in2(_gnd_net_),
            .in3(N__20717),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_22_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_22_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_22_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_22_3  (
            .in0(N__20691),
            .in1(N__20636),
            .in2(_gnd_net_),
            .in3(N__20603),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_22_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21059),
            .in3(N__21023),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_22_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_22_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_22_5  (
            .in0(_gnd_net_),
            .in1(N__21016),
            .in2(_gnd_net_),
            .in3(N__20984),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_22_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_22_6  (
            .in0(_gnd_net_),
            .in1(N__20977),
            .in2(_gnd_net_),
            .in3(N__20948),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_22_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(N__20944),
            .in2(_gnd_net_),
            .in3(N__20915),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_23_0  (
            .in0(_gnd_net_),
            .in1(N__21159),
            .in2(_gnd_net_),
            .in3(N__20903),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(N__21081),
            .in2(_gnd_net_),
            .in3(N__20885),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(N__21120),
            .in2(_gnd_net_),
            .in3(N__20873),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20870),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_23_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_23_4  (
            .in0(_gnd_net_),
            .in1(N__21160),
            .in2(_gnd_net_),
            .in3(N__21175),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_23_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_23_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_23_5  (
            .in0(N__21121),
            .in1(_gnd_net_),
            .in2(N__21145),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_6  (
            .in0(N__22588),
            .in1(N__22558),
            .in2(_gnd_net_),
            .in3(N__26027),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_23_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_23_7  (
            .in0(_gnd_net_),
            .in1(N__21082),
            .in2(_gnd_net_),
            .in3(N__21097),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un7_start_stop_LC_2_30_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.un7_start_stop_LC_2_30_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un7_start_stop_LC_2_30_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.un7_start_stop_LC_2_30_3  (
            .in0(N__30007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49269),
            .lcout(un7_start_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_1 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_1  (
            .in0(N__23270),
            .in1(N__25479),
            .in2(N__23474),
            .in3(N__22232),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50033),
            .ce(),
            .sr(N__49204));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_3_12_2  (
            .in0(N__21989),
            .in1(N__23453),
            .in2(_gnd_net_),
            .in3(N__23272),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50033),
            .ce(),
            .sr(N__49204));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_12_7 .LUT_INIT=16'b0011001011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_3_12_7  (
            .in0(N__23271),
            .in1(N__22039),
            .in2(N__23475),
            .in3(N__23660),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50033),
            .ce(),
            .sr(N__49204));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_13_0 .LUT_INIT=16'b1100110011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_3_13_0  (
            .in0(N__25512),
            .in1(N__22094),
            .in2(N__23476),
            .in3(N__23274),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50022),
            .ce(),
            .sr(N__49208));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_13_5 .LUT_INIT=16'b1011000010110001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_3_13_5  (
            .in0(N__23273),
            .in1(N__25514),
            .in2(N__22208),
            .in3(N__23466),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50022),
            .ce(),
            .sr(N__49208));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_3_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_3_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_3_13_6 .LUT_INIT=16'b1100110001000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_3_13_6  (
            .in0(N__25513),
            .in1(N__21887),
            .in2(N__23477),
            .in3(N__23275),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50022),
            .ce(),
            .sr(N__49208));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_1 .LUT_INIT=16'b1111001111100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_1  (
            .in0(N__23436),
            .in1(N__23264),
            .in2(N__22073),
            .in3(N__25522),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50011),
            .ce(),
            .sr(N__49212));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_3_14_6 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_3_14_6  (
            .in0(N__25521),
            .in1(N__23437),
            .in2(N__23285),
            .in3(N__22298),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50011),
            .ce(),
            .sr(N__49212));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_3_15_2 .LUT_INIT=16'b1101110011011000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_3_15_2  (
            .in0(N__23258),
            .in1(N__21968),
            .in2(N__25523),
            .in3(N__23423),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50000),
            .ce(),
            .sr(N__49217));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_3 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_3  (
            .in0(N__23420),
            .in1(N__25516),
            .in2(N__22289),
            .in3(N__23262),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50000),
            .ce(),
            .sr(N__49217));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_4 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_4  (
            .in0(N__25515),
            .in1(N__23422),
            .in2(N__23284),
            .in3(N__22271),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50000),
            .ce(),
            .sr(N__49217));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_5 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_5  (
            .in0(N__23421),
            .in1(N__25517),
            .in2(N__22262),
            .in3(N__23263),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50000),
            .ce(),
            .sr(N__49217));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__21218),
            .in2(N__21254),
            .in3(N__21242),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__21545),
            .in2(N__21212),
            .in3(N__21200),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__21500),
            .in2(N__21536),
            .in3(N__21524),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_16_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_16_3  (
            .in0(N__21494),
            .in1(N__21458),
            .in2(N__21470),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_16_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_16_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_16_4  (
            .in0(N__21452),
            .in1(N__21419),
            .in2(N__21428),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_16_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(N__21377),
            .in2(N__21413),
            .in3(N__21401),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_16_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(N__21338),
            .in2(N__21371),
            .in3(N__21362),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_16_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_16_7  (
            .in0(_gnd_net_),
            .in1(N__21299),
            .in2(N__21332),
            .in3(N__21323),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__21260),
            .in2(N__21293),
            .in3(N__21284),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__21629),
            .in2(N__21662),
            .in3(N__21653),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_3_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_3_17_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_3_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21623),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49979),
            .ce(),
            .sr(N__49228));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_18_1  (
            .in0(N__23848),
            .in1(N__23932),
            .in2(N__24028),
            .in3(N__23796),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_18_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_18_2  (
            .in0(N__24115),
            .in1(N__24197),
            .in2(N__21596),
            .in3(N__24276),
            .lcout(\current_shift_inst.PI_CTRL.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_3_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_3_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_3_19_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_3_19_0  (
            .in0(N__30421),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49964),
            .ce(),
            .sr(N__49237));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30199),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49964),
            .ce(),
            .sr(N__49237));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30133),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49964),
            .ce(),
            .sr(N__49237));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30481),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49964),
            .ce(),
            .sr(N__49237));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_20_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_20_7 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_20_7  (
            .in0(N__21793),
            .in1(N__21745),
            .in2(N__21719),
            .in3(N__21866),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_21_0  (
            .in0(N__22508),
            .in1(N__22625),
            .in2(N__22502),
            .in3(N__22514),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ),
            .ltout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_21_1 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__25235),
            .in2(N__21689),
            .in3(N__21674),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_21_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(N__23973),
            .in2(_gnd_net_),
            .in3(N__25180),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_21_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(N__25179),
            .in2(_gnd_net_),
            .in3(N__24066),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_21_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_21_5  (
            .in0(N__23974),
            .in1(N__25353),
            .in2(N__21686),
            .in3(N__23901),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(\current_shift_inst.PI_CTRL.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_21_6 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_21_6  (
            .in0(N__25236),
            .in1(N__24157),
            .in2(N__21683),
            .in3(N__25269),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_0  (
            .in0(N__23902),
            .in1(N__21680),
            .in2(N__24071),
            .in3(N__25354),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_3_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_3_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_3_22_1 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_3_22_1  (
            .in0(N__25268),
            .in1(N__24156),
            .in2(N__25240),
            .in3(N__21673),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_22_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_22_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_22_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_22_2  (
            .in0(_gnd_net_),
            .in1(N__22056),
            .in2(_gnd_net_),
            .in3(N__21708),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_22_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_22_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_22_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_22_3  (
            .in0(N__25317),
            .in1(N__21837),
            .in2(N__21878),
            .in3(N__25108),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_22_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_3_22_4  (
            .in0(N__25109),
            .in1(N__25318),
            .in2(N__21844),
            .in3(N__22057),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_22_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_22_5  (
            .in0(_gnd_net_),
            .in1(N__24155),
            .in2(_gnd_net_),
            .in3(N__24237),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_22_6 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_22_6  (
            .in0(N__21808),
            .in1(N__25227),
            .in2(N__21857),
            .in3(N__25139),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(\current_shift_inst.PI_CTRL.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_3_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_3_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_3_22_7 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_3_22_7  (
            .in0(N__21763),
            .in1(N__21854),
            .in2(N__21848),
            .in3(N__24238),
            .lcout(\current_shift_inst.PI_CTRL.N_160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_3_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_3_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_3_23_0 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_3_23_0  (
            .in0(N__25241),
            .in1(N__23975),
            .in2(N__25152),
            .in3(N__25281),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(),
            .sr(N__49246));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_3_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_3_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_3_23_1 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_3_23_1  (
            .in0(N__24158),
            .in1(N__21821),
            .in2(N__21812),
            .in3(N__25147),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(),
            .sr(N__49246));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_3_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_3_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_3_23_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_3_23_4  (
            .in0(N__24239),
            .in1(N__21764),
            .in2(_gnd_net_),
            .in3(N__21752),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(),
            .sr(N__49246));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_3_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_3_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_3_23_5 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_3_23_5  (
            .in0(N__25280),
            .in1(N__25243),
            .in2(N__25154),
            .in3(N__24070),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(),
            .sr(N__49246));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_3_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_3_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_3_23_6 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_3_23_6  (
            .in0(N__25242),
            .in1(N__23903),
            .in2(N__25153),
            .in3(N__25282),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(),
            .sr(N__49246));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_4_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_4_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_4_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29126),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50046),
            .ce(),
            .sr(N__49183));
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_4_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_4_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__23651),
            .in2(N__22040),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__22019),
            .in2(N__23613),
            .in3(N__22007),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__24255),
            .in2(N__22004),
            .in3(N__21983),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__21980),
            .in2(N__24208),
            .in3(N__21956),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__24111),
            .in2(N__21953),
            .in3(N__21923),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(N__24003),
            .in2(N__21920),
            .in3(N__21905),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(N__23921),
            .in2(N__21902),
            .in3(N__21881),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__23834),
            .in2(N__22250),
            .in3(N__22226),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__23789),
            .in2(N__22223),
            .in3(N__22199),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__23736),
            .in2(N__22196),
            .in3(N__22181),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__24733),
            .in2(N__22178),
            .in3(N__22145),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__22142),
            .in2(N__24668),
            .in3(N__22130),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__24614),
            .in2(N__22127),
            .in3(N__22112),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(N__24551),
            .in2(N__22109),
            .in3(N__22088),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__22085),
            .in2(N__24500),
            .in3(N__22064),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__24446),
            .in2(N__22784),
            .in3(N__22304),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__24396),
            .in2(N__22733),
            .in3(N__22301),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__24329),
            .in2(N__22682),
            .in3(N__22292),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__22637),
            .in2(N__25065),
            .in3(N__22280),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__25010),
            .in2(N__23093),
            .in3(N__22277),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__24962),
            .in2(N__23057),
            .in3(N__22274),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(N__24911),
            .in2(N__23021),
            .in3(N__22265),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(N__22988),
            .in2(N__24865),
            .in3(N__22253),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(N__24814),
            .in2(N__22955),
            .in3(N__22352),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__25877),
            .in2(N__22922),
            .in3(N__22349),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__22886),
            .in2(N__25996),
            .in3(N__22346),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__25953),
            .in2(N__22862),
            .in3(N__22343),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__25914),
            .in2(N__23576),
            .in3(N__22340),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__25617),
            .in2(N__23540),
            .in3(N__22337),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__25563),
            .in2(N__23507),
            .in3(N__22334),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_15_6  (
            .in0(N__27032),
            .in1(N__25408),
            .in2(N__23492),
            .in3(N__22331),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_16_0 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_4_16_0  (
            .in0(N__23425),
            .in1(N__25505),
            .in2(N__22328),
            .in3(N__23181),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(),
            .sr(N__49218));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_4_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_4_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_4_16_1 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_4_16_1  (
            .in0(N__25503),
            .in1(N__23429),
            .in2(N__23222),
            .in3(N__22439),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(),
            .sr(N__49218));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_4_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_4_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_4_16_2 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_4_16_2  (
            .in0(N__23424),
            .in1(N__25507),
            .in2(N__22433),
            .in3(N__23168),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(),
            .sr(N__49218));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_4_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_4_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_4_16_3 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_4_16_3  (
            .in0(N__25501),
            .in1(N__23427),
            .in2(N__23220),
            .in3(N__22421),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(),
            .sr(N__49218));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_4 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_4  (
            .in0(N__23426),
            .in1(N__25506),
            .in2(N__22415),
            .in3(N__23182),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(),
            .sr(N__49218));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_4_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_4_16_5 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_4_16_5  (
            .in0(N__25504),
            .in1(N__23430),
            .in2(N__23223),
            .in3(N__22406),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(),
            .sr(N__49218));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_4_16_7 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_4_16_7  (
            .in0(N__25502),
            .in1(N__23428),
            .in2(N__23221),
            .in3(N__22400),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49980),
            .ce(),
            .sr(N__49218));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_17_0  (
            .in0(N__22379),
            .in1(N__22358),
            .in2(N__22394),
            .in3(N__22478),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_17_2  (
            .in0(N__25616),
            .in1(N__24628),
            .in2(N__24508),
            .in3(N__23757),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_17_3 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_17_3  (
            .in0(N__23806),
            .in1(N__22472),
            .in2(N__22373),
            .in3(N__24029),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_17_6  (
            .in0(N__25064),
            .in1(N__24916),
            .in2(N__24400),
            .in3(N__24333),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_17_7  (
            .in0(N__25404),
            .in1(N__24864),
            .in2(N__22481),
            .in3(N__23702),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_18_0 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_18_0  (
            .in0(N__24277),
            .in1(N__23623),
            .in2(N__24207),
            .in3(N__23673),
            .lcout(\current_shift_inst.PI_CTRL.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1  (
            .in0(N__24501),
            .in1(N__24627),
            .in2(N__23761),
            .in3(N__24454),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_2  (
            .in0(N__24679),
            .in1(N__22466),
            .in2(N__22457),
            .in3(N__25567),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_18_4  (
            .in0(N__24915),
            .in1(N__24337),
            .in2(N__25069),
            .in3(N__24392),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_18_5  (
            .in0(N__25618),
            .in1(N__24863),
            .in2(N__22454),
            .in3(N__22451),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_19_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(N__23690),
            .in2(_gnd_net_),
            .in3(N__23674),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49955),
            .ce(),
            .sr(N__49234));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_20_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_20_1  (
            .in0(N__23723),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24640),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_20_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_20_2  (
            .in0(N__25643),
            .in1(N__24695),
            .in2(N__22442),
            .in3(N__22619),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_20_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_20_3  (
            .in0(N__24418),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24469),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_20_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_20_5  (
            .in0(N__23722),
            .in1(N__25592),
            .in2(N__24419),
            .in3(N__24470),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_20_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_20_6  (
            .in0(N__24641),
            .in1(N__24694),
            .in2(N__22517),
            .in3(N__22493),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_21_0  (
            .in0(N__24833),
            .in1(N__24787),
            .in2(N__24593),
            .in3(N__24526),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_21_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_21_1  (
            .in0(N__24772),
            .in1(N__24985),
            .in2(N__24757),
            .in3(N__25030),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_21_2  (
            .in0(N__25031),
            .in1(N__24527),
            .in2(N__24989),
            .in3(N__24592),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_21_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_21_3  (
            .in0(_gnd_net_),
            .in1(N__24304),
            .in2(_gnd_net_),
            .in3(N__24358),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_21_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_21_4  (
            .in0(N__24887),
            .in1(N__24773),
            .in2(N__24761),
            .in3(N__22487),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_21_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_21_5  (
            .in0(_gnd_net_),
            .in1(N__24886),
            .in2(_gnd_net_),
            .in3(N__24937),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_21_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_21_6  (
            .in0(N__25661),
            .in1(N__25639),
            .in2(N__22628),
            .in3(N__25537),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_21_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_21_7  (
            .in0(N__25588),
            .in1(N__24832),
            .in2(N__24788),
            .in3(N__24938),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_22_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_22_6  (
            .in0(N__25660),
            .in1(N__24305),
            .in2(N__24362),
            .in3(N__25538),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_22_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_22_7  (
            .in0(N__22613),
            .in1(N__22604),
            .in2(N__22598),
            .in3(N__22595),
            .lcout(\current_shift_inst.PI_CTRL.N_158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_4_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_4_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_4_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_4_23_6  (
            .in0(_gnd_net_),
            .in1(N__25082),
            .in2(_gnd_net_),
            .in3(N__26040),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49244));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_4_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_4_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_4_23_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_4_23_7  (
            .in0(N__26041),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22568),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49244));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_5_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_5_12_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_5_12_7  (
            .in0(N__22538),
            .in1(N__23438),
            .in2(_gnd_net_),
            .in3(N__23268),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50012),
            .ce(),
            .sr(N__49194));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_5_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_5_13_1 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_5_13_1  (
            .in0(N__23281),
            .in1(N__25475),
            .in2(N__23473),
            .in3(N__22532),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50001),
            .ce(),
            .sr(N__49200));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_5_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_5_13_2 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_5_13_2  (
            .in0(N__25471),
            .in1(N__23440),
            .in2(N__22526),
            .in3(N__23283),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50001),
            .ce(),
            .sr(N__49200));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_5_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_5_13_3 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_5_13_3  (
            .in0(N__23278),
            .in1(N__25472),
            .in2(N__23470),
            .in3(N__22850),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50001),
            .ce(),
            .sr(N__49200));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_5_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_5_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_5_13_5 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_5_13_5  (
            .in0(N__23280),
            .in1(N__25474),
            .in2(N__23472),
            .in3(N__22844),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50001),
            .ce(),
            .sr(N__49200));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_13_6 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_5_13_6  (
            .in0(N__25470),
            .in1(N__23439),
            .in2(N__22838),
            .in3(N__23282),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50001),
            .ce(),
            .sr(N__49200));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_13_7 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_5_13_7  (
            .in0(N__23279),
            .in1(N__25473),
            .in2(N__23471),
            .in3(N__22829),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50001),
            .ce(),
            .sr(N__49200));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_5_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_5_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__22823),
            .in2(N__22808),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_5_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_5_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__22772),
            .in2(N__22751),
            .in3(N__22724),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_5_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_5_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__22721),
            .in2(N__22700),
            .in3(N__22673),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_5_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_5_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__22670),
            .in2(N__22652),
            .in3(N__22631),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_5_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_5_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__23108),
            .in2(N__27110),
            .in3(N__23081),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_5_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_5_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__23078),
            .in2(N__27112),
            .in3(N__23045),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_5_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_5_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__23042),
            .in2(N__27111),
            .in3(N__23012),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_5_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_5_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__23009),
            .in2(N__27113),
            .in3(N__22982),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_5_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_5_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__27090),
            .in2(N__22979),
            .in3(N__22946),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_5_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_5_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__22943),
            .in2(N__27114),
            .in3(N__22913),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_5_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__27094),
            .in2(N__22910),
            .in3(N__22880),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_5_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_5_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__22877),
            .in2(N__27115),
            .in3(N__22853),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_5_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_5_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__23591),
            .in2(N__27120),
            .in3(N__23564),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_5_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_5_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(N__23561),
            .in2(N__27116),
            .in3(N__23531),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_5_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_5_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(N__23528),
            .in2(N__27121),
            .in3(N__23498),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_5_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_5_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23495),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_5_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_5_16_2 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_5_16_2  (
            .in0(N__23385),
            .in1(N__25435),
            .in2(N__23224),
            .in3(N__23483),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49970),
            .ce(),
            .sr(N__49213));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_4 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_4  (
            .in0(N__23386),
            .in1(N__25436),
            .in2(N__23225),
            .in3(N__23309),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49970),
            .ce(),
            .sr(N__49213));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_17_0  (
            .in0(N__23696),
            .in1(N__23303),
            .in2(N__25850),
            .in3(N__23291),
            .lcout(\current_shift_inst.PI_CTRL.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_17_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_17_1  (
            .in0(N__25910),
            .in1(N__25949),
            .in2(N__25881),
            .in3(N__25559),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_5_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_5_17_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(N__25985),
            .in2(_gnd_net_),
            .in3(N__24963),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_5_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_5_17_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_5_17_6  (
            .in0(N__24806),
            .in1(N__25011),
            .in2(N__23711),
            .in3(N__23708),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_17_7  (
            .in0(N__25012),
            .in1(N__24807),
            .in2(N__24974),
            .in3(N__25403),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30166),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(),
            .sr(N__49223));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30106),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(),
            .sr(N__49223));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30452),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(),
            .sr(N__49223));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30070),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(),
            .sr(N__49223));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__23689),
            .in2(N__23675),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__23630),
            .in2(N__23624),
            .in3(N__23594),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49229));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__24290),
            .in2(N__24281),
            .in3(N__24218),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49229));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_19_3  (
            .in0(_gnd_net_),
            .in1(N__24215),
            .in2(N__24209),
            .in3(N__24125),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49229));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_19_4  (
            .in0(_gnd_net_),
            .in1(N__24122),
            .in2(N__24116),
            .in3(N__24032),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49229));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_19_5  (
            .in0(_gnd_net_),
            .in1(N__24024),
            .in2(N__23987),
            .in3(N__23948),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49229));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(N__23945),
            .in2(N__23939),
            .in3(N__23867),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49229));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_19_7  (
            .in0(_gnd_net_),
            .in1(N__23864),
            .in2(N__23855),
            .in3(N__23813),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49229));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(N__25802),
            .in2(N__23810),
            .in3(N__23765),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__49941),
            .ce(),
            .sr(N__49235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_20_1  (
            .in0(_gnd_net_),
            .in1(N__26273),
            .in2(N__23762),
            .in3(N__23714),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__49941),
            .ce(),
            .sr(N__49235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_20_2  (
            .in0(_gnd_net_),
            .in1(N__25823),
            .in2(N__24740),
            .in3(N__24686),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__49941),
            .ce(),
            .sr(N__49235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_20_3  (
            .in0(_gnd_net_),
            .in1(N__26264),
            .in2(N__24683),
            .in3(N__24632),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__49941),
            .ce(),
            .sr(N__49235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_20_4  (
            .in0(_gnd_net_),
            .in1(N__25814),
            .in2(N__24629),
            .in3(N__24578),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__49941),
            .ce(),
            .sr(N__49235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_20_5  (
            .in0(_gnd_net_),
            .in1(N__26282),
            .in2(N__24575),
            .in3(N__24518),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__49941),
            .ce(),
            .sr(N__49235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_20_6  (
            .in0(_gnd_net_),
            .in1(N__27020),
            .in2(N__24515),
            .in3(N__24461),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__49941),
            .ce(),
            .sr(N__49235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_20_7  (
            .in0(_gnd_net_),
            .in1(N__24458),
            .in2(N__27839),
            .in3(N__24407),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__49941),
            .ce(),
            .sr(N__49235));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_21_0  (
            .in0(_gnd_net_),
            .in1(N__26246),
            .in2(N__24404),
            .in3(N__24347),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_5_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49238));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_21_1  (
            .in0(_gnd_net_),
            .in1(N__26993),
            .in2(N__24344),
            .in3(N__24293),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49238));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_21_2  (
            .in0(_gnd_net_),
            .in1(N__26255),
            .in2(N__25076),
            .in3(N__25022),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49238));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_21_3  (
            .in0(_gnd_net_),
            .in1(N__27011),
            .in2(N__25019),
            .in3(N__24977),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49238));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_21_4  (
            .in0(_gnd_net_),
            .in1(N__27002),
            .in2(N__24973),
            .in3(N__24929),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49238));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_21_5  (
            .in0(_gnd_net_),
            .in1(N__27827),
            .in2(N__24926),
            .in3(N__24878),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49238));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_21_6  (
            .in0(_gnd_net_),
            .in1(N__26237),
            .in2(N__24875),
            .in3(N__24824),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49238));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_21_7  (
            .in0(_gnd_net_),
            .in1(N__29057),
            .in2(N__24821),
            .in3(N__24776),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49238));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_22_0  (
            .in0(_gnd_net_),
            .in1(N__27947),
            .in2(N__25889),
            .in3(N__24764),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_5_22_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49239));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_22_1  (
            .in0(_gnd_net_),
            .in1(N__27818),
            .in2(N__26000),
            .in3(N__25664),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49239));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_22_2  (
            .in0(_gnd_net_),
            .in1(N__26984),
            .in2(N__25964),
            .in3(N__25646),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49239));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(N__29030),
            .in2(N__25928),
            .in3(N__25628),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49239));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_22_4  (
            .in0(_gnd_net_),
            .in1(N__29048),
            .in2(N__25625),
            .in3(N__25577),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49239));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_22_5  (
            .in0(_gnd_net_),
            .in1(N__29039),
            .in2(N__25574),
            .in3(N__25526),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__49929),
            .ce(),
            .sr(N__49239));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_22_6  (
            .in0(N__27956),
            .in1(N__25511),
            .in2(_gnd_net_),
            .in3(N__25358),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49929),
            .ce(),
            .sr(N__49239));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_5_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_5_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_5_23_0 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_5_23_0  (
            .in0(N__25214),
            .in1(N__25140),
            .in2(N__25355),
            .in3(N__25288),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49923),
            .ce(),
            .sr(N__49240));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_5_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_5_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_5_23_1 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_5_23_1  (
            .in0(N__25289),
            .in1(N__25215),
            .in2(N__25181),
            .in3(N__25151),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49923),
            .ce(),
            .sr(N__49240));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25835),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49923),
            .ce(),
            .sr(N__49240));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_9_2 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_7_9_2  (
            .in0(N__28820),
            .in1(N__25708),
            .in2(_gnd_net_),
            .in3(N__29118),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_LC_7_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_7_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_7_9_3 .LUT_INIT=16'b1000101011111010;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_7_9_3  (
            .in0(N__25709),
            .in1(N__28747),
            .in2(N__25712),
            .in3(N__28821),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50023),
            .ce(),
            .sr(N__49168));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__28766),
            .in2(_gnd_net_),
            .in3(N__26221),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_9_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__28819),
            .in2(_gnd_net_),
            .in3(N__28743),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_9_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25700),
            .in3(N__28767),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__26456),
            .in2(N__25697),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_7_10_1  (
            .in0(N__26196),
            .in1(N__26414),
            .in2(_gnd_net_),
            .in3(N__25685),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__50013),
            .ce(),
            .sr(N__49173));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_7_10_2  (
            .in0(N__26204),
            .in1(N__26381),
            .in2(N__25682),
            .in3(N__25670),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__50013),
            .ce(),
            .sr(N__49173));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_10_3  (
            .in0(N__26197),
            .in1(N__26348),
            .in2(_gnd_net_),
            .in3(N__25667),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__50013),
            .ce(),
            .sr(N__49173));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_7_10_4  (
            .in0(N__26205),
            .in1(N__26672),
            .in2(_gnd_net_),
            .in3(N__25739),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__50013),
            .ce(),
            .sr(N__49173));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_7_10_5  (
            .in0(N__26198),
            .in1(N__26651),
            .in2(_gnd_net_),
            .in3(N__25736),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__50013),
            .ce(),
            .sr(N__49173));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_7_10_6  (
            .in0(N__26206),
            .in1(N__26618),
            .in2(_gnd_net_),
            .in3(N__25733),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__50013),
            .ce(),
            .sr(N__49173));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_7_10_7  (
            .in0(N__26199),
            .in1(N__26597),
            .in2(_gnd_net_),
            .in3(N__25730),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__50013),
            .ce(),
            .sr(N__49173));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_7_11_0  (
            .in0(N__26203),
            .in1(N__26570),
            .in2(_gnd_net_),
            .in3(N__25727),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__50002),
            .ce(),
            .sr(N__49179));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_7_11_1  (
            .in0(N__26192),
            .in1(N__26537),
            .in2(_gnd_net_),
            .in3(N__25724),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__50002),
            .ce(),
            .sr(N__49179));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_7_11_2  (
            .in0(N__26200),
            .in1(N__26519),
            .in2(_gnd_net_),
            .in3(N__25721),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__50002),
            .ce(),
            .sr(N__49179));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_7_11_3  (
            .in0(N__26193),
            .in1(N__26489),
            .in2(_gnd_net_),
            .in3(N__25718),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__50002),
            .ce(),
            .sr(N__49179));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_7_11_4  (
            .in0(N__26201),
            .in1(N__26768),
            .in2(_gnd_net_),
            .in3(N__25715),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__50002),
            .ce(),
            .sr(N__49179));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_7_11_5  (
            .in0(N__26194),
            .in1(N__26749),
            .in2(_gnd_net_),
            .in3(N__25766),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__50002),
            .ce(),
            .sr(N__49179));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_7_11_6  (
            .in0(N__26202),
            .in1(N__26723),
            .in2(_gnd_net_),
            .in3(N__25763),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__50002),
            .ce(),
            .sr(N__49179));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_7  (
            .in0(N__26195),
            .in1(N__27211),
            .in2(_gnd_net_),
            .in3(N__25760),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__50002),
            .ce(),
            .sr(N__49179));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_7_12_0  (
            .in0(N__26173),
            .in1(N__27238),
            .in2(_gnd_net_),
            .in3(N__25757),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49989),
            .ce(),
            .sr(N__49184));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_7_12_1  (
            .in0(N__26177),
            .in1(N__26298),
            .in2(_gnd_net_),
            .in3(N__25754),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49989),
            .ce(),
            .sr(N__49184));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_7_12_2  (
            .in0(N__26174),
            .in1(N__26319),
            .in2(_gnd_net_),
            .in3(N__25751),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49989),
            .ce(),
            .sr(N__49184));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_7_12_3  (
            .in0(N__26178),
            .in1(N__26842),
            .in2(_gnd_net_),
            .in3(N__25748),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49989),
            .ce(),
            .sr(N__49184));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_7_12_4  (
            .in0(N__26175),
            .in1(N__26824),
            .in2(_gnd_net_),
            .in3(N__25745),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49989),
            .ce(),
            .sr(N__49184));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_7_12_5  (
            .in0(N__26179),
            .in1(N__27321),
            .in2(_gnd_net_),
            .in3(N__25742),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49989),
            .ce(),
            .sr(N__49184));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_7_12_6  (
            .in0(N__26176),
            .in1(N__27295),
            .in2(_gnd_net_),
            .in3(N__25793),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49989),
            .ce(),
            .sr(N__49184));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_7_12_7  (
            .in0(N__26180),
            .in1(N__27744),
            .in2(_gnd_net_),
            .in3(N__25790),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49989),
            .ce(),
            .sr(N__49184));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_7_13_0  (
            .in0(N__26169),
            .in1(N__27777),
            .in2(_gnd_net_),
            .in3(N__25787),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49981),
            .ce(),
            .sr(N__49189));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_7_13_1  (
            .in0(N__26207),
            .in1(N__26930),
            .in2(_gnd_net_),
            .in3(N__25784),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49981),
            .ce(),
            .sr(N__49189));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_7_13_2  (
            .in0(N__26170),
            .in1(N__26947),
            .in2(_gnd_net_),
            .in3(N__25781),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49981),
            .ce(),
            .sr(N__49189));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_7_13_3  (
            .in0(N__26208),
            .in1(N__27565),
            .in2(_gnd_net_),
            .in3(N__25778),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49981),
            .ce(),
            .sr(N__49189));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_7_13_4  (
            .in0(N__26171),
            .in1(N__27594),
            .in2(_gnd_net_),
            .in3(N__25775),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49981),
            .ce(),
            .sr(N__49189));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_7_13_5  (
            .in0(N__26209),
            .in1(N__27489),
            .in2(_gnd_net_),
            .in3(N__25772),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49981),
            .ce(),
            .sr(N__49189));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_7_13_6  (
            .in0(N__26172),
            .in1(N__27519),
            .in2(_gnd_net_),
            .in3(N__25769),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49981),
            .ce(),
            .sr(N__49189));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_14_0 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_14_0  (
            .in0(N__31235),
            .in1(N__31196),
            .in2(N__31167),
            .in3(N__32688),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49971),
            .ce(),
            .sr(N__49195));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_7_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_7_14_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__31954),
            .in2(_gnd_net_),
            .in3(N__38392),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_14_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26003),
            .in3(N__36696),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__28834),
            .in2(_gnd_net_),
            .in3(N__29119),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_7_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_7_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_7_16_3  (
            .in0(N__25995),
            .in1(N__25957),
            .in2(N__25924),
            .in3(N__25882),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29632),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49936),
            .ce(),
            .sr(N__49219));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30322),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(),
            .sr(N__49224));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30268),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(),
            .sr(N__49224));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_20_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_7_20_4  (
            .in0(N__30379),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(),
            .sr(N__49224));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30235),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(),
            .sr(N__49224));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30352),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(),
            .sr(N__49224));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_20_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(N__30298),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(),
            .sr(N__49224));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_7_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_7_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30592),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49924),
            .ce(),
            .sr(N__49230));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30655),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49924),
            .ce(),
            .sr(N__49230));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_7_21_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_7_21_5  (
            .in0(N__30967),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49924),
            .ce(),
            .sr(N__49230));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_7_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_7_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_7_22_2  (
            .in0(_gnd_net_),
            .in1(N__36700),
            .in2(_gnd_net_),
            .in3(N__36724),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_22_3 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_7_22_3  (
            .in0(N__28783),
            .in1(N__26228),
            .in2(N__26443),
            .in3(N__26181),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(),
            .sr(N__49236));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_7_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_7_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_7_22_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_7_22_6  (
            .in0(_gnd_net_),
            .in1(N__26057),
            .in2(_gnd_net_),
            .in3(N__26045),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(),
            .sr(N__49236));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_8_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_8_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_8_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_8_6_4  (
            .in0(N__35370),
            .in1(N__28393),
            .in2(_gnd_net_),
            .in3(N__32411),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50040),
            .ce(N__28913),
            .sr(N__49146));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_8_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_8_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_8_7_3  (
            .in0(N__32357),
            .in1(N__29180),
            .in2(_gnd_net_),
            .in3(N__33838),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50034),
            .ce(N__28914),
            .sr(N__49153));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_8_8_0  (
            .in0(N__27188),
            .in1(N__34469),
            .in2(_gnd_net_),
            .in3(N__32330),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50024),
            .ce(N__28915),
            .sr(N__49158));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_8_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_8_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_8_8_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_8_8_1  (
            .in0(N__32328),
            .in1(N__28044),
            .in2(N__34400),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50024),
            .ce(N__28915),
            .sr(N__49158));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_8_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_8_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_8_8_2  (
            .in0(N__28506),
            .in1(N__33617),
            .in2(_gnd_net_),
            .in3(N__32332),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50024),
            .ce(N__28915),
            .sr(N__49158));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_8_8_4  (
            .in0(N__33476),
            .in1(N__27173),
            .in2(_gnd_net_),
            .in3(N__32333),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50024),
            .ce(N__28915),
            .sr(N__49158));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_8_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_8_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_8_8_5  (
            .in0(N__32329),
            .in1(N__27270),
            .in2(_gnd_net_),
            .in3(N__35015),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50024),
            .ce(N__28915),
            .sr(N__49158));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_8_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_8_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_8_8_6  (
            .in0(N__29417),
            .in1(N__34646),
            .in2(_gnd_net_),
            .in3(N__32331),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50024),
            .ce(N__28915),
            .sr(N__49158));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_8_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_8_9_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_8_9_0  (
            .in0(N__26321),
            .in1(N__26299),
            .in2(N__26468),
            .in3(N__26330),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_8_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_8_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_8_9_1  (
            .in0(N__26329),
            .in1(N__26320),
            .in2(N__26303),
            .in3(N__26464),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_8_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_8_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_8_9_3  (
            .in0(N__31076),
            .in1(N__34942),
            .in2(_gnd_net_),
            .in3(N__32405),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50014),
            .ce(N__28916),
            .sr(N__49163));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_8_9_4  (
            .in0(N__32404),
            .in1(N__29204),
            .in2(_gnd_net_),
            .in3(N__29240),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50014),
            .ce(N__28916),
            .sr(N__49163));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_8_9_5  (
            .in0(N__27988),
            .in1(N__33908),
            .in2(_gnd_net_),
            .in3(N__32406),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50014),
            .ce(N__28916),
            .sr(N__49163));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_8_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_8_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_8_9_7  (
            .in0(N__33768),
            .in1(N__28589),
            .in2(_gnd_net_),
            .in3(N__32407),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50014),
            .ce(N__28916),
            .sr(N__49163));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_8_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_8_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__27374),
            .in2(N__26423),
            .in3(N__26455),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_8_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_8_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_8_10_1  (
            .in0(N__26413),
            .in1(N__26402),
            .in2(N__26396),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_8_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_8_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__26387),
            .in2(N__26369),
            .in3(N__26380),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_8_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_8_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__26336),
            .in2(N__26360),
            .in3(N__26347),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_8_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_8_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__26678),
            .in2(N__26660),
            .in3(N__26671),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_8_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_8_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__26777),
            .in2(N__26639),
            .in3(N__26650),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_8_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_8_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__26627),
            .in2(N__26606),
            .in3(N__26617),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_8_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_8_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__26585),
            .in2(N__26972),
            .in3(N__26596),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_8_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_8_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__26579),
            .in2(N__26558),
            .in3(N__26569),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_8_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_8_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__26525),
            .in2(N__26549),
            .in3(N__26536),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_8_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_8_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_8_11_2  (
            .in0(N__26518),
            .in1(N__26507),
            .in2(N__26498),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_8_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_8_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__27644),
            .in2(N__26477),
            .in3(N__26488),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_8_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_8_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__26756),
            .in2(N__27431),
            .in3(N__26767),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_8_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_8_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__27422),
            .in2(N__26735),
            .in3(N__26750),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_8_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_8_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__26711),
            .in2(N__27404),
            .in3(N__26722),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_8_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_8_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__27251),
            .in2(N__27197),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_8_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_8_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__26705),
            .in2(N__26693),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_8_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_8_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__26852),
            .in2(N__26807),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_8_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_8_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__27281),
            .in2(N__27368),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_8_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_8_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__27158),
            .in2(N__27722),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_8_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_8_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__26915),
            .in2(N__26960),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_8_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_8_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__27530),
            .in2(N__26885),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_8_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_8_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__27470),
            .in2(N__26870),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26855),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_13_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_8_13_0  (
            .in0(N__26786),
            .in1(N__26795),
            .in2(N__26843),
            .in3(N__26823),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_13_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_8_13_1  (
            .in0(N__26794),
            .in1(N__26841),
            .in2(N__26825),
            .in3(N__26785),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_8_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_8_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_8_13_2  (
            .in0(N__32359),
            .in1(N__27889),
            .in2(_gnd_net_),
            .in3(N__34852),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49972),
            .ce(N__28919),
            .sr(N__49185));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_8_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_8_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_8_13_3  (
            .in0(N__34784),
            .in1(N__31310),
            .in2(_gnd_net_),
            .in3(N__32362),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49972),
            .ce(N__28919),
            .sr(N__49185));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_8_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_8_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_8_13_4  (
            .in0(N__32360),
            .in1(N__28638),
            .in2(_gnd_net_),
            .in3(N__33689),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49972),
            .ce(N__28919),
            .sr(N__49185));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_8_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_8_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_8_13_5  (
            .in0(N__33544),
            .in1(N__28471),
            .in2(_gnd_net_),
            .in3(N__32358),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(elapsed_time_ns_1_RNIKJ91B_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_8_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_8_13_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_8_13_6  (
            .in0(N__32361),
            .in1(_gnd_net_),
            .in2(N__26975),
            .in3(N__33545),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49972),
            .ce(N__28919),
            .sr(N__49185));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_14_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_14_0  (
            .in0(N__26929),
            .in1(N__26906),
            .in2(N__26897),
            .in3(N__26946),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_14_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_8_14_1  (
            .in0(N__26905),
            .in1(N__26896),
            .in2(N__26948),
            .in3(N__26928),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_8_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_8_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_8_14_2  (
            .in0(N__27860),
            .in1(N__35531),
            .in2(_gnd_net_),
            .in3(N__32421),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49965),
            .ce(N__28921),
            .sr(N__49190));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_8_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_8_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_8_14_3  (
            .in0(N__32419),
            .in1(N__35441),
            .in2(_gnd_net_),
            .in3(N__27464),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49965),
            .ce(N__28921),
            .sr(N__49190));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_8_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_8_14_6 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_8_14_6  (
            .in0(N__27623),
            .in1(N__27564),
            .in2(N__27598),
            .in3(N__27544),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_8_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_8_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_8_14_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_8_14_7  (
            .in0(N__32420),
            .in1(N__35276),
            .in2(_gnd_net_),
            .in3(N__28427),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49965),
            .ce(N__28921),
            .sr(N__49190));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_15_4 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_8_15_4  (
            .in0(N__27679),
            .in1(N__27520),
            .in2(N__27496),
            .in3(N__27694),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_16_0 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_8_16_0  (
            .in0(N__27709),
            .in1(N__27784),
            .in2(N__27757),
            .in3(N__28937),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_8_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_8_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__27146),
            .in2(_gnd_net_),
            .in3(N__27125),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_8_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_8_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_8_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30721),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49925),
            .ce(),
            .sr(N__49220));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_8_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_8_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_8_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30565),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49917),
            .ce(),
            .sr(N__49225));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_8_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_8_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30535),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49917),
            .ce(),
            .sr(N__49225));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_8_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_8_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_8_21_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_8_21_6  (
            .in0(_gnd_net_),
            .in1(N__30622),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49917),
            .ce(),
            .sr(N__49225));
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_8_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_8_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_8_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_27_LC_8_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30844),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49231));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_9_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_9_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_9_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_9_5_4  (
            .in0(N__27275),
            .in1(N__35014),
            .in2(_gnd_net_),
            .in3(N__32410),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50041),
            .ce(N__32737),
            .sr(N__49135));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_2  (
            .in0(N__34718),
            .in1(N__28027),
            .in2(_gnd_net_),
            .in3(N__32409),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50035),
            .ce(N__28912),
            .sr(N__49139));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_7_2  (
            .in0(N__32353),
            .in1(N__34467),
            .in2(_gnd_net_),
            .in3(N__27187),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_7_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_9_7_3  (
            .in0(N__34468),
            .in1(_gnd_net_),
            .in2(N__27176),
            .in3(N__32355),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50025),
            .ce(N__32738),
            .sr(N__49147));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_9_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_9_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_9_7_5  (
            .in0(N__33474),
            .in1(N__27172),
            .in2(_gnd_net_),
            .in3(N__32352),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(elapsed_time_ns_1_RNILK91B_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_7_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_9_7_6  (
            .in0(N__32354),
            .in1(_gnd_net_),
            .in2(N__27161),
            .in3(N__33475),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50025),
            .ce(N__32738),
            .sr(N__49147));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_7_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_9_7_7  (
            .in0(N__27660),
            .in1(_gnd_net_),
            .in2(N__34319),
            .in3(N__32356),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50025),
            .ce(N__32738),
            .sr(N__49147));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_8_0  (
            .in0(N__32304),
            .in1(N__27664),
            .in2(_gnd_net_),
            .in3(N__34315),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_8_1  (
            .in0(N__29271),
            .in1(N__27394),
            .in2(_gnd_net_),
            .in3(N__32307),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_8_2  (
            .in0(N__32306),
            .in1(N__28507),
            .in2(_gnd_net_),
            .in3(N__33616),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_8_3  (
            .in0(N__27989),
            .in1(N__33903),
            .in2(_gnd_net_),
            .in3(N__32308),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_4  (
            .in0(N__33902),
            .in1(N__29239),
            .in2(N__33839),
            .in3(N__29270),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_9_8_5  (
            .in0(N__31309),
            .in1(N__34776),
            .in2(_gnd_net_),
            .in3(N__32303),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_9_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_9_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_9_8_6  (
            .in0(N__32309),
            .in1(N__28046),
            .in2(_gnd_net_),
            .in3(N__34396),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_8_7  (
            .in0(N__27274),
            .in1(N__35007),
            .in2(_gnd_net_),
            .in3(N__32305),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_9_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_9_9_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_9_9_2  (
            .in0(N__32397),
            .in1(_gnd_net_),
            .in2(N__27890),
            .in3(N__34856),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50003),
            .ce(N__32721),
            .sr(N__49159));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_9_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_9_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_9_9_3  (
            .in0(N__34101),
            .in1(N__27415),
            .in2(_gnd_net_),
            .in3(N__32394),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(elapsed_time_ns_1_RNI2COBB_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_9_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_9_9_4  (
            .in0(N__32395),
            .in1(_gnd_net_),
            .in2(N__27254),
            .in3(N__34102),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50003),
            .ce(N__32721),
            .sr(N__49159));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_9_5 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_9_5  (
            .in0(N__27634),
            .in1(N__31871),
            .in2(N__31285),
            .in3(N__31901),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6  (
            .in0(N__32396),
            .in1(N__27390),
            .in2(_gnd_net_),
            .in3(N__29272),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50003),
            .ce(N__32721),
            .sr(N__49159));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_9_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_9_10_0 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_9_10_0  (
            .in0(N__27452),
            .in1(N__27220),
            .in2(N__27443),
            .in3(N__27245),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_9_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_9_10_1 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_9_10_1  (
            .in0(N__27244),
            .in1(N__27451),
            .in2(N__27224),
            .in3(N__27439),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_9_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_9_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_9_10_2  (
            .in0(N__32400),
            .in1(N__29348),
            .in2(_gnd_net_),
            .in3(N__34044),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49990),
            .ce(N__28917),
            .sr(N__49164));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_9_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_9_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_9_10_3  (
            .in0(N__33974),
            .in1(N__32401),
            .in2(_gnd_net_),
            .in3(N__29381),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49990),
            .ce(N__28917),
            .sr(N__49164));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_9_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_9_10_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_9_10_4  (
            .in0(N__32398),
            .in1(_gnd_net_),
            .in2(N__29315),
            .in3(N__34244),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49990),
            .ce(N__28917),
            .sr(N__49164));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_9_10_5  (
            .in0(N__32006),
            .in1(N__34174),
            .in2(_gnd_net_),
            .in3(N__32402),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49990),
            .ce(N__28917),
            .sr(N__49164));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_9_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_9_10_6  (
            .in0(N__32399),
            .in1(N__34106),
            .in2(_gnd_net_),
            .in3(N__27416),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49990),
            .ce(N__28917),
            .sr(N__49164));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_9_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_9_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_9_10_7  (
            .in0(N__29273),
            .in1(N__27395),
            .in2(_gnd_net_),
            .in3(N__32403),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49990),
            .ce(N__28917),
            .sr(N__49164));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_11_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_9_11_0  (
            .in0(N__27328),
            .in1(N__27347),
            .in2(N__27305),
            .in3(N__27359),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_11_1 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_9_11_1  (
            .in0(N__27358),
            .in1(N__27346),
            .in2(N__27332),
            .in3(N__27304),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_9_11_7  (
            .in0(N__27668),
            .in1(N__34304),
            .in2(_gnd_net_),
            .in3(N__32408),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49982),
            .ce(N__28918),
            .sr(N__49169));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0  (
            .in0(N__27638),
            .in1(N__31870),
            .in2(N__31286),
            .in3(N__31900),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_12_1  (
            .in0(N__32393),
            .in1(N__33687),
            .in2(_gnd_net_),
            .in3(N__28639),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_9_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_9_12_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_9_12_2  (
            .in0(N__29307),
            .in1(N__32392),
            .in2(_gnd_net_),
            .in3(N__34239),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_5 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_9_12_5  (
            .in0(N__27622),
            .in1(N__27599),
            .in2(N__27572),
            .in3(N__27545),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_12_6 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_9_12_6  (
            .in0(N__27524),
            .in1(N__27683),
            .in2(N__27500),
            .in3(N__27698),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_13_0 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_9_13_0  (
            .in0(N__31712),
            .in1(N__27794),
            .in2(N__27806),
            .in3(N__31732),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_9_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_9_13_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_9_13_1  (
            .in0(N__27793),
            .in1(N__31711),
            .in2(N__31736),
            .in3(N__27802),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_13_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_13_2  (
            .in0(N__35429),
            .in1(N__32417),
            .in2(_gnd_net_),
            .in3(N__27463),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_9_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_9_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_9_13_3 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_9_13_3  (
            .in0(N__32418),
            .in1(N__35430),
            .in2(N__27809),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49966),
            .ce(N__32679),
            .sr(N__49180));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_9_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_9_13_7 .LUT_INIT=16'b1000101011101111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_9_13_7  (
            .in0(N__32473),
            .in1(N__28666),
            .in2(N__32771),
            .in3(N__28654),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_9_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_9_14_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_9_14_1  (
            .in0(N__27859),
            .in1(N__35525),
            .in2(_gnd_net_),
            .in3(N__32426),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49957),
            .ce(N__32560),
            .sr(N__49186));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_9_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_9_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_9_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_9_14_5  (
            .in0(N__32449),
            .in1(N__34577),
            .in2(_gnd_net_),
            .in3(N__32425),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49957),
            .ce(N__32560),
            .sr(N__49186));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_15_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_15_0  (
            .in0(N__27710),
            .in1(N__27785),
            .in2(N__27758),
            .in3(N__28936),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_15_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_9_15_2  (
            .in0(N__32453),
            .in1(N__32423),
            .in2(_gnd_net_),
            .in3(N__34576),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49948),
            .ce(N__28922),
            .sr(N__49191));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_15_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_9_15_4  (
            .in0(N__35149),
            .in1(N__32424),
            .in2(_gnd_net_),
            .in3(N__28975),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49948),
            .ce(N__28922),
            .sr(N__49191));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_9_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_9_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_9_15_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_9_15_7  (
            .in0(N__32422),
            .in1(N__28561),
            .in2(_gnd_net_),
            .in3(N__35192),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49948),
            .ce(N__28922),
            .sr(N__49191));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_9_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_9_16_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__29807),
            .in2(_gnd_net_),
            .in3(N__31945),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_9_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_9_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_9_16_1  (
            .in0(N__27882),
            .in1(N__34845),
            .in2(_gnd_net_),
            .in3(N__32415),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_9_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_9_16_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_9_16_7  (
            .in0(N__27858),
            .in1(N__35527),
            .in2(_gnd_net_),
            .in3(N__32416),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_17_0 .LUT_INIT=16'b1000101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_9_17_0  (
            .in0(N__31946),
            .in1(N__28866),
            .in2(N__38399),
            .in3(N__36692),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49201));
    defparam \phase_controller_inst2.start_timer_hc_LC_9_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_9_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_9_17_1 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_9_17_1  (
            .in0(N__28847),
            .in1(N__28678),
            .in2(N__29813),
            .in3(N__33353),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49201));
    defparam \phase_controller_inst2.state_2_LC_9_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_9_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_9_17_2 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst2.state_2_LC_9_17_2  (
            .in0(N__29934),
            .in1(N__28883),
            .in2(N__29891),
            .in3(N__28867),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49201));
    defparam \phase_controller_inst1.state_4_LC_9_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_9_17_3 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_9_17_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_9_17_3  (
            .in0(N__29995),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33352),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49201));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29808),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49201));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_9_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_9_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_9_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30691),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49214));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_9_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_9_21_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__30508),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49913),
            .ce(),
            .sr(N__49221));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_9_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_9_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_9_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30871),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49909),
            .ce(),
            .sr(N__49226));
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_31_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30737),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49909),
            .ce(),
            .sr(N__49226));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_9_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_9_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_9_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30901),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49909),
            .ce(),
            .sr(N__49226));
    defparam \phase_controller_inst2.S1_LC_9_28_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_28_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_28_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29887),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49895),
            .ce(),
            .sr(N__49245));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_6 (
            .in0(N__27929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_10_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_10_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_10_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_10_5_3  (
            .in0(N__31072),
            .in1(N__34943),
            .in2(_gnd_net_),
            .in3(N__32327),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50027),
            .ce(N__32736),
            .sr(N__49122));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_6_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_6_0  (
            .in0(N__31534),
            .in1(N__27911),
            .in2(N__27902),
            .in3(N__31507),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_6_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_10_6_1  (
            .in0(N__27910),
            .in1(N__31535),
            .in2(N__31508),
            .in3(N__27901),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_6_2  (
            .in0(N__32325),
            .in1(N__35374),
            .in2(_gnd_net_),
            .in3(N__28392),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_6_7  (
            .in0(N__28028),
            .in1(N__34716),
            .in2(_gnd_net_),
            .in3(N__32326),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_10_7_0  (
            .in0(N__34645),
            .in1(N__29412),
            .in2(_gnd_net_),
            .in3(N__32186),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__32702),
            .sr(N__49136));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_10_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_10_7_2  (
            .in0(N__28045),
            .in1(N__34395),
            .in2(_gnd_net_),
            .in3(N__32185),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__32702),
            .sr(N__49136));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_10_7_3  (
            .in0(N__32184),
            .in1(N__28026),
            .in2(_gnd_net_),
            .in3(N__34717),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__32702),
            .sr(N__49136));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_10_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_10_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_10_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_10_7_4  (
            .in0(N__29196),
            .in1(N__29229),
            .in2(_gnd_net_),
            .in3(N__32187),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__32702),
            .sr(N__49136));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_10_7_6  (
            .in0(N__29175),
            .in1(N__33834),
            .in2(_gnd_net_),
            .in3(N__32188),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50004),
            .ce(N__32702),
            .sr(N__49136));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0  (
            .in0(N__31843),
            .in1(N__28001),
            .in2(N__31819),
            .in3(N__28010),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1  (
            .in0(N__28009),
            .in1(N__28000),
            .in2(N__31820),
            .in3(N__31844),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_10_8_6  (
            .in0(N__27987),
            .in1(N__33907),
            .in2(_gnd_net_),
            .in3(N__32190),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49992),
            .ce(N__32726),
            .sr(N__49140));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_10_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_10_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__27962),
            .in2(N__27971),
            .in3(N__31172),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_10_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_10_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__28160),
            .in2(N__28151),
            .in3(N__31127),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_10_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_10_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__28142),
            .in2(N__28136),
            .in3(N__31100),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_10_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_10_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__28127),
            .in2(N__28118),
            .in3(N__31478),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_10_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_10_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__28607),
            .in2(N__28109),
            .in3(N__31457),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_10_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_10_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_10_9_5  (
            .in0(N__31436),
            .in1(N__28100),
            .in2(N__28619),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_10_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_10_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__28487),
            .in2(N__28094),
            .in3(N__31415),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_10_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_10_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__28460),
            .in2(N__28085),
            .in3(N__31394),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_10_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_10_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__28073),
            .in2(N__28064),
            .in3(N__31373),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_10_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_10_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__28055),
            .in2(N__28283),
            .in3(N__31352),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_10_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_10_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__28274),
            .in2(N__28262),
            .in3(N__31331),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_10_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_10_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__28253),
            .in2(N__28241),
            .in3(N__31667),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_10_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_10_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__29288),
            .in2(N__28232),
            .in3(N__31646),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_10_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_10_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__28598),
            .in2(N__28223),
            .in3(N__31625),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_10_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_10_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__28205),
            .in2(N__28214),
            .in3(N__31604),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_10_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_10_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__29396),
            .in2(N__29390),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_10_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_10_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__28199),
            .in2(N__28190),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_10_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_10_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__28178),
            .in2(N__28172),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_10_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_10_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__28352),
            .in2(N__28343),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_10_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_10_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__28289),
            .in2(N__28520),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_10_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_10_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__28328),
            .in2(N__28319),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_10_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_10_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__28436),
            .in2(N__28448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_10_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_10_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__28361),
            .in2(N__28307),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28292),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_12_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_10_12_0  (
            .in0(N__28544),
            .in1(N__31760),
            .in2(N__31787),
            .in3(N__28529),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_10_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_10_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_10_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_10_12_3  (
            .in0(N__28958),
            .in1(N__34508),
            .in2(_gnd_net_),
            .in3(N__32345),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49959),
            .ce(N__32687),
            .sr(N__49165));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_12_4 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_10_12_4  (
            .in0(N__28543),
            .in1(N__31759),
            .in2(N__31786),
            .in3(N__28528),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_10_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_10_12_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_10_12_6  (
            .in0(N__32344),
            .in1(N__33609),
            .in2(_gnd_net_),
            .in3(N__28511),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49959),
            .ce(N__32687),
            .sr(N__49165));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_10_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_10_12_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_10_12_7  (
            .in0(N__33538),
            .in1(N__28478),
            .in2(_gnd_net_),
            .in3(N__32346),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49959),
            .ce(N__32687),
            .sr(N__49165));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_13_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_13_0  (
            .in0(N__32792),
            .in1(N__31687),
            .in2(N__28406),
            .in3(N__28370),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_13_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_13_1  (
            .in0(N__28369),
            .in1(N__32791),
            .in2(N__31691),
            .in3(N__28402),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_13_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_13_2  (
            .in0(N__35270),
            .in1(N__32338),
            .in2(_gnd_net_),
            .in3(N__28420),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(elapsed_time_ns_1_RNI7IPBB_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_10_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_10_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_10_13_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_10_13_3  (
            .in0(N__32340),
            .in1(_gnd_net_),
            .in2(N__28409),
            .in3(N__35271),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49950),
            .ce(N__32631),
            .sr(N__49170));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_13_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_10_13_5  (
            .in0(N__32339),
            .in1(N__35363),
            .in2(_gnd_net_),
            .in3(N__28394),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49950),
            .ce(N__32631),
            .sr(N__49170));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_13_7 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_13_7  (
            .in0(N__32474),
            .in1(N__28667),
            .in2(N__32770),
            .in3(N__28655),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_10_14_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_10_14_2  (
            .in0(N__32347),
            .in1(N__28560),
            .in2(_gnd_net_),
            .in3(N__35191),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__32627),
            .sr(N__49174));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_10_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_10_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_10_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_10_14_4  (
            .in0(N__32348),
            .in1(N__35148),
            .in2(_gnd_net_),
            .in3(N__28974),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__32627),
            .sr(N__49174));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_10_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_10_14_5  (
            .in0(N__33688),
            .in1(N__28643),
            .in2(_gnd_net_),
            .in3(N__32351),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__32627),
            .sr(N__49174));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_10_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_10_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_10_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_10_14_6  (
            .in0(N__32349),
            .in1(N__33770),
            .in2(_gnd_net_),
            .in3(N__28578),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__32627),
            .sr(N__49174));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_10_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_10_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_10_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_10_14_7  (
            .in0(N__32002),
            .in1(N__34175),
            .in2(_gnd_net_),
            .in3(N__32350),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__32627),
            .sr(N__49174));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_15_0  (
            .in0(N__32335),
            .in1(N__28957),
            .in2(_gnd_net_),
            .in3(N__34513),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_2  (
            .in0(N__32334),
            .in1(N__33769),
            .in2(_gnd_net_),
            .in3(N__28582),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_10_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_10_15_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__29584),
            .in2(_gnd_net_),
            .in3(N__29462),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_15_5  (
            .in0(N__28562),
            .in1(N__35190),
            .in2(_gnd_net_),
            .in3(N__32336),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_15_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_10_15_7  (
            .in0(N__28976),
            .in1(N__35147),
            .in2(_gnd_net_),
            .in3(N__32337),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_10_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_10_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_10_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_10_16_1  (
            .in0(N__28953),
            .in1(N__34514),
            .in2(_gnd_net_),
            .in3(N__32414),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49931),
            .ce(N__28920),
            .sr(N__49187));
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_10_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_10_17_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_RNIG7JF_2_LC_10_17_2  (
            .in0(N__28882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28862),
            .lcout(\phase_controller_inst2.N_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_17_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_10_17_3  (
            .in0(N__28702),
            .in1(N__28881),
            .in2(N__28868),
            .in3(N__29015),
            .lcout(\phase_controller_inst2.N_51_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__29785),
            .in2(_gnd_net_),
            .in3(N__35994),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_165_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_10_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_10_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__29935),
            .in2(_gnd_net_),
            .in3(N__29874),
            .lcout(\phase_controller_inst2.test_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_10_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_10_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_10_18_0 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst2.state_0_LC_10_18_0  (
            .in0(N__29086),
            .in1(N__28711),
            .in2(N__29072),
            .in3(N__29020),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49920),
            .ce(),
            .sr(N__49196));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_10_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_10_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_10_18_3 .LUT_INIT=16'b1000110010101100;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_10_18_3  (
            .in0(N__28841),
            .in1(N__29087),
            .in2(N__28790),
            .in3(N__28748),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49920),
            .ce(),
            .sr(N__49196));
    defparam \phase_controller_inst2.state_1_LC_10_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_10_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_10_18_5 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.state_1_LC_10_18_5  (
            .in0(N__28712),
            .in1(N__29019),
            .in2(_gnd_net_),
            .in3(N__28679),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49920),
            .ce(),
            .sr(N__49196));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_18_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_18_6 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_10_18_6  (
            .in0(N__29786),
            .in1(N__35966),
            .in2(_gnd_net_),
            .in3(N__35996),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49920),
            .ce(),
            .sr(N__49196));
    defparam \phase_controller_inst2.start_timer_tr_LC_10_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_10_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_10_18_7 .LUT_INIT=16'b0011001101110011;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_10_18_7  (
            .in0(N__33351),
            .in1(N__29132),
            .in2(N__29117),
            .in3(N__29902),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49920),
            .ce(),
            .sr(N__49196));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_10_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_10_19_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__29085),
            .in2(_gnd_net_),
            .in3(N__29068),
            .lcout(\phase_controller_inst2.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_10_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_10_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_10_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30928),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49906),
            .ce(),
            .sr(N__49209));
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_10_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_10_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_10_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_29_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30784),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49215));
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_10_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_10_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_10_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_30_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30757),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49215));
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_10_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_10_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_10_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_28_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30808),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49215));
    defparam \phase_controller_inst2.S2_LC_10_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_10_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_10_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29021),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49900),
            .ce(),
            .sr(N__49222));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_6_5 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_6_5  (
            .in0(N__31022),
            .in1(N__33207),
            .in2(N__31049),
            .in3(N__35814),
            .lcout(\phase_controller_inst1.N_49_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33934),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49993),
            .ce(N__35099),
            .sr(N__49129));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33865),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49993),
            .ce(N__35099),
            .sr(N__49129));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_11_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_11_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_11_7_5  (
            .in0(N__29200),
            .in1(N__29228),
            .in2(_gnd_net_),
            .in3(N__32165),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_11_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_11_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_11_7_7  (
            .in0(N__29179),
            .in1(N__33830),
            .in2(_gnd_net_),
            .in3(N__32166),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_11_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_11_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_11_8_0  (
            .in0(N__34385),
            .in1(N__34458),
            .in2(N__34314),
            .in3(N__33465),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_11_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_11_8_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__33537),
            .in2(_gnd_net_),
            .in3(N__33608),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_11_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_11_8_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_11_8_2  (
            .in0(N__33683),
            .in1(N__33758),
            .in2(N__29159),
            .in3(N__29156),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_11_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_11_8_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_11_8_4  (
            .in0(N__35375),
            .in1(N__35440),
            .in2(_gnd_net_),
            .in3(N__29150),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_11_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_11_8_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_11_8_5  (
            .in0(N__35150),
            .in1(N__29141),
            .in2(N__29135),
            .in3(N__30977),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_8_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_11_8_6  (
            .in0(N__29416),
            .in1(_gnd_net_),
            .in2(N__29420),
            .in3(N__34640),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_8_7  (
            .in0(N__29344),
            .in1(N__34045),
            .in2(_gnd_net_),
            .in3(N__32164),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_11_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_11_9_0 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_11_9_0  (
            .in0(N__29324),
            .in1(N__31579),
            .in2(N__29360),
            .in3(N__31556),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_11_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_11_9_1 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_11_9_1  (
            .in0(N__31555),
            .in1(N__29323),
            .in2(N__31583),
            .in3(N__29356),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_11_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_11_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_11_9_2  (
            .in0(N__33969),
            .in1(N__32167),
            .in2(_gnd_net_),
            .in3(N__29374),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(elapsed_time_ns_1_RNI4EOBB_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_11_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_11_9_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_11_9_3  (
            .in0(N__32169),
            .in1(_gnd_net_),
            .in2(N__29363),
            .in3(N__33970),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49974),
            .ce(N__32703),
            .sr(N__49141));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_11_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_11_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_11_9_5  (
            .in0(N__32168),
            .in1(N__29340),
            .in2(_gnd_net_),
            .in3(N__34046),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49974),
            .ce(N__32703),
            .sr(N__49141));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_11_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_11_9_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_11_9_6  (
            .in0(N__29314),
            .in1(N__32170),
            .in2(_gnd_net_),
            .in3(N__34243),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49974),
            .ce(N__32703),
            .sr(N__49141));
    defparam \phase_controller_inst1.start_timer_tr_LC_11_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_11_10_1 .LUT_INIT=16'b0101010101011101;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_11_10_1  (
            .in0(N__29282),
            .in1(N__29454),
            .in2(N__33374),
            .in3(N__31979),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49967),
            .ce(),
            .sr(N__49148));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_10_2 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_10_2  (
            .in0(N__29453),
            .in1(N__29470),
            .in2(_gnd_net_),
            .in3(N__29571),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_LC_11_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_11_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_11_10_3 .LUT_INIT=16'b1011101000111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_11_10_3  (
            .in0(N__29471),
            .in1(N__29577),
            .in2(N__29474),
            .in3(N__29548),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49967),
            .ce(),
            .sr(N__49148));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_11_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_11_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_11_10_4  (
            .in0(N__29455),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49967),
            .ce(),
            .sr(N__49148));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_11_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_11_10_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__29570),
            .in2(_gnd_net_),
            .in3(N__29544),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_11_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_11_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29438),
            .in3(N__31218),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_11_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_11_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_11_11_0  (
            .in0(N__29749),
            .in1(N__33927),
            .in2(_gnd_net_),
            .in3(N__29435),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__49960),
            .ce(N__29857),
            .sr(N__49154));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_11_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_11_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_11_11_1  (
            .in0(N__29745),
            .in1(N__33864),
            .in2(_gnd_net_),
            .in3(N__29432),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__49960),
            .ce(N__29857),
            .sr(N__49154));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_11_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_11_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_11_11_2  (
            .in0(N__29750),
            .in1(N__33784),
            .in2(_gnd_net_),
            .in3(N__29429),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__49960),
            .ce(N__29857),
            .sr(N__49154));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_11_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_11_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_11_11_3  (
            .in0(N__29746),
            .in1(N__33705),
            .in2(_gnd_net_),
            .in3(N__29426),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__49960),
            .ce(N__29857),
            .sr(N__49154));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_11_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_11_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_11_11_4  (
            .in0(N__29751),
            .in1(N__33633),
            .in2(_gnd_net_),
            .in3(N__29423),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__49960),
            .ce(N__29857),
            .sr(N__49154));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_11_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_11_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_11_11_5  (
            .in0(N__29747),
            .in1(N__33561),
            .in2(_gnd_net_),
            .in3(N__29501),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__49960),
            .ce(N__29857),
            .sr(N__49154));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_11_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_11_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_11_11_6  (
            .in0(N__29752),
            .in1(N__33490),
            .in2(_gnd_net_),
            .in3(N__29498),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__49960),
            .ce(N__29857),
            .sr(N__49154));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_11_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_11_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_11_11_7  (
            .in0(N__29748),
            .in1(N__33417),
            .in2(_gnd_net_),
            .in3(N__29495),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__49960),
            .ce(N__29857),
            .sr(N__49154));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_11_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_11_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_11_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_11_12_0  (
            .in0(N__29709),
            .in1(N__34428),
            .in2(_gnd_net_),
            .in3(N__29492),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__49951),
            .ce(N__29858),
            .sr(N__49160));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_11_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_11_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_11_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_11_12_1  (
            .in0(N__29738),
            .in1(N__34347),
            .in2(_gnd_net_),
            .in3(N__29489),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__49951),
            .ce(N__29858),
            .sr(N__49160));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_11_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_11_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_11_12_2  (
            .in0(N__29706),
            .in1(N__34260),
            .in2(_gnd_net_),
            .in3(N__29486),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__49951),
            .ce(N__29858),
            .sr(N__49160));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_11_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_11_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_11_12_3  (
            .in0(N__29735),
            .in1(N__34191),
            .in2(_gnd_net_),
            .in3(N__29483),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__49951),
            .ce(N__29858),
            .sr(N__49160));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_11_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_11_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_11_12_4  (
            .in0(N__29707),
            .in1(N__34122),
            .in2(_gnd_net_),
            .in3(N__29480),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__49951),
            .ce(N__29858),
            .sr(N__49160));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_11_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_11_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_11_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_11_12_5  (
            .in0(N__29736),
            .in1(N__34062),
            .in2(_gnd_net_),
            .in3(N__29477),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__49951),
            .ce(N__29858),
            .sr(N__49160));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_11_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_11_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_11_12_6  (
            .in0(N__29708),
            .in1(N__33990),
            .in2(_gnd_net_),
            .in3(N__29528),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__49951),
            .ce(N__29858),
            .sr(N__49160));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_11_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_11_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_11_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_11_12_7  (
            .in0(N__29737),
            .in1(N__35029),
            .in2(_gnd_net_),
            .in3(N__29525),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__49951),
            .ce(N__29858),
            .sr(N__49160));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_11_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_11_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_11_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_11_13_0  (
            .in0(N__29731),
            .in1(N__34965),
            .in2(_gnd_net_),
            .in3(N__29522),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__49944),
            .ce(N__29856),
            .sr(N__49166));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_11_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_11_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_11_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_11_13_1  (
            .in0(N__29762),
            .in1(N__34878),
            .in2(_gnd_net_),
            .in3(N__29519),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__49944),
            .ce(N__29856),
            .sr(N__49166));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_11_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_11_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_11_13_2  (
            .in0(N__29732),
            .in1(N__34800),
            .in2(_gnd_net_),
            .in3(N__29516),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__49944),
            .ce(N__29856),
            .sr(N__49166));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_11_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_11_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_11_13_3  (
            .in0(N__29763),
            .in1(N__34734),
            .in2(_gnd_net_),
            .in3(N__29513),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__49944),
            .ce(N__29856),
            .sr(N__49166));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_11_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_11_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_11_13_4  (
            .in0(N__29733),
            .in1(N__34662),
            .in2(_gnd_net_),
            .in3(N__29510),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__49944),
            .ce(N__29856),
            .sr(N__49166));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_11_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_11_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_11_13_5  (
            .in0(N__29764),
            .in1(N__34591),
            .in2(_gnd_net_),
            .in3(N__29507),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__49944),
            .ce(N__29856),
            .sr(N__49166));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_11_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_11_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_11_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_11_13_6  (
            .in0(N__29734),
            .in1(N__34528),
            .in2(_gnd_net_),
            .in3(N__29504),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__49944),
            .ce(N__29856),
            .sr(N__49166));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_11_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_11_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_11_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_11_13_7  (
            .in0(N__29765),
            .in1(N__35545),
            .in2(_gnd_net_),
            .in3(N__29606),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__49944),
            .ce(N__29856),
            .sr(N__49166));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_11_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_11_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_11_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_11_14_0  (
            .in0(N__29739),
            .in1(N__35463),
            .in2(_gnd_net_),
            .in3(N__29603),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__49939),
            .ce(N__29852),
            .sr(N__49171));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_11_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_11_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_11_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_11_14_1  (
            .in0(N__29743),
            .in1(N__35391),
            .in2(_gnd_net_),
            .in3(N__29600),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__49939),
            .ce(N__29852),
            .sr(N__49171));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_11_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_11_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_11_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_11_14_2  (
            .in0(N__29740),
            .in1(N__35292),
            .in2(_gnd_net_),
            .in3(N__29597),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__49939),
            .ce(N__29852),
            .sr(N__49171));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_11_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_11_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_11_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_11_14_3  (
            .in0(N__29744),
            .in1(N__35206),
            .in2(_gnd_net_),
            .in3(N__29594),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__49939),
            .ce(N__29852),
            .sr(N__49171));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_11_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_11_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_11_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_11_14_4  (
            .in0(N__29741),
            .in1(N__35317),
            .in2(_gnd_net_),
            .in3(N__29591),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__49939),
            .ce(N__29852),
            .sr(N__49171));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_11_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_11_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_11_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_11_14_5  (
            .in0(N__35233),
            .in1(N__29742),
            .in2(_gnd_net_),
            .in3(N__29588),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49939),
            .ce(N__29852),
            .sr(N__49171));
    defparam \phase_controller_inst1.state_0_LC_11_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_11_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_11_15_1 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_0_LC_11_15_1  (
            .in0(N__33211),
            .in1(N__30020),
            .in2(N__30038),
            .in3(N__35825),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(),
            .sr(N__49175));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_11_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_11_15_2 .LUT_INIT=16'b1000110010101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_11_15_2  (
            .in0(N__29585),
            .in1(N__30037),
            .in2(N__31234),
            .in3(N__29552),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(),
            .sr(N__49175));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__30033),
            .in2(_gnd_net_),
            .in3(N__30019),
            .lcout(\phase_controller_inst1.N_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNILR64_4_LC_11_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNILR64_4_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNILR64_4_LC_11_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNILR64_4_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__29994),
            .in2(_gnd_net_),
            .in3(N__33363),
            .lcout(phase_controller_inst1_N_54),
            .ltout(phase_controller_inst1_N_54_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_3_LC_11_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_11_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_11_16_6 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst2.state_3_LC_11_16_6  (
            .in0(N__29880),
            .in1(N__29942),
            .in2(N__29909),
            .in3(N__29906),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(),
            .sr(N__49181));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_17_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_17_0  (
            .in0(N__29784),
            .in1(N__35965),
            .in2(_gnd_net_),
            .in3(N__35995),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_17_2 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_17_2  (
            .in0(N__29812),
            .in1(N__31912),
            .in2(_gnd_net_),
            .in3(N__31950),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_11_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_11_17_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_11_17_4  (
            .in0(N__29783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_11_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_11_18_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_11_18_0  (
            .in0(N__37016),
            .in1(N__38579),
            .in2(_gnd_net_),
            .in3(N__41802),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_11_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_11_18_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_11_18_2  (
            .in0(N__38516),
            .in1(N__36953),
            .in2(_gnd_net_),
            .in3(N__41800),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_18_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29639),
            .in3(N__32935),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(),
            .sr(N__49192));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41801),
            .lcout(\current_shift_inst.N_1271_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_11_18_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_11_18_7  (
            .in0(N__41803),
            .in1(N__38564),
            .in2(_gnd_net_),
            .in3(N__37001),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_11_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_11_19_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_11_19_0  (
            .in0(N__32915),
            .in1(N__30212),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_11_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_11_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_11_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__32906),
            .in2(_gnd_net_),
            .in3(N__30173),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49197));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_11_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_11_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_11_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32894),
            .in3(N__30140),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49197));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_11_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_11_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_11_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__32879),
            .in2(_gnd_net_),
            .in3(N__30110),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49197));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_11_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_11_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_11_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__32867),
            .in2(_gnd_net_),
            .in3(N__30074),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49197));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_11_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_11_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_11_19_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32855),
            .in3(N__30041),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49197));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_11_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_11_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_11_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__32840),
            .in2(_gnd_net_),
            .in3(N__30455),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49197));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_11_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_11_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_11_19_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32828),
            .in3(N__30425),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49197));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_11_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_11_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_11_20_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32807),
            .in3(N__30392),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__49907),
            .ce(),
            .sr(N__49202));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_11_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_11_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_11_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__33056),
            .in2(_gnd_net_),
            .in3(N__30362),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__49907),
            .ce(),
            .sr(N__49202));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_11_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_11_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_11_20_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33044),
            .in3(N__30332),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__49907),
            .ce(),
            .sr(N__49202));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_11_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_11_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_11_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__33029),
            .in2(_gnd_net_),
            .in3(N__30302),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__49907),
            .ce(),
            .sr(N__49202));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_11_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_11_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_11_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(N__33017),
            .in2(_gnd_net_),
            .in3(N__30278),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__49907),
            .ce(),
            .sr(N__49202));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_11_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_11_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_11_20_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33005),
            .in3(N__30245),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__49907),
            .ce(),
            .sr(N__49202));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_11_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_11_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_11_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__32990),
            .in2(_gnd_net_),
            .in3(N__30215),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__49907),
            .ce(),
            .sr(N__49202));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_11_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_11_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_11_20_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32978),
            .in3(N__30701),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__49907),
            .ce(),
            .sr(N__49202));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_11_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_11_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_11_21_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32963),
            .in3(N__30665),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__49904),
            .ce(),
            .sr(N__49205));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_11_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_11_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_11_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__33173),
            .in2(_gnd_net_),
            .in3(N__30635),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__49904),
            .ce(),
            .sr(N__49205));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_11_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_11_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_11_21_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33161),
            .in3(N__30602),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__49904),
            .ce(),
            .sr(N__49205));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_11_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_11_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_11_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__33146),
            .in2(_gnd_net_),
            .in3(N__30572),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__49904),
            .ce(),
            .sr(N__49205));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_11_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_11_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_11_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__33134),
            .in2(_gnd_net_),
            .in3(N__30545),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__49904),
            .ce(),
            .sr(N__49205));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_11_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_11_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_11_21_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33122),
            .in3(N__30515),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__49904),
            .ce(),
            .sr(N__49205));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_11_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_11_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_11_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__33107),
            .in2(_gnd_net_),
            .in3(N__30491),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__49904),
            .ce(),
            .sr(N__49205));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_11_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_11_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_11_21_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33095),
            .in3(N__30944),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__49904),
            .ce(),
            .sr(N__49205));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_11_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_11_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_11_22_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33080),
            .in3(N__30914),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49210));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_11_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_11_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_11_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__33314),
            .in2(_gnd_net_),
            .in3(N__30884),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49210));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_11_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_11_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_11_22_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33302),
            .in3(N__30851),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49210));
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_11_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_11_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_11_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_27_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__33287),
            .in2(_gnd_net_),
            .in3(N__30824),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49210));
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_11_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_11_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_11_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_28_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__33275),
            .in2(_gnd_net_),
            .in3(N__30794),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49210));
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_11_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_11_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_11_22_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_29_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33263),
            .in3(N__30767),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49210));
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_11_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_11_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_11_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_30_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__33230),
            .in2(_gnd_net_),
            .in3(N__30743),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ),
            .clk(N__49901),
            .ce(),
            .sr(N__49210));
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_11_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_11_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_11_22_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_31_LC_11_22_7  (
            .in0(N__33245),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30740),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49901),
            .ce(),
            .sr(N__49210));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_12_3_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_12_3_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_12_3_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_12_3_2  (
            .in0(N__44305),
            .in1(N__44276),
            .in2(_gnd_net_),
            .in3(N__50527),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50026),
            .ce(N__49521),
            .sr(N__49099));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_12_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_12_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_12_5_2  (
            .in0(N__50484),
            .in1(N__40248),
            .in2(_gnd_net_),
            .in3(N__43368),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_12_5_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_12_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_12_5_4  (
            .in0(N__31071),
            .in1(N__34935),
            .in2(_gnd_net_),
            .in3(N__32324),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_12_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_12_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_12_6_0 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_2_LC_12_6_0  (
            .in0(N__31047),
            .in1(N__35667),
            .in2(N__31028),
            .in3(N__35886),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49991),
            .ce(),
            .sr(N__49115));
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_12_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_12_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNIE87F_2_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__31023),
            .in2(_gnd_net_),
            .in3(N__31046),
            .lcout(\phase_controller_inst1.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_3 .LUT_INIT=16'b1000110010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_3  (
            .in0(N__39551),
            .in1(N__31048),
            .in2(N__39455),
            .in3(N__39504),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49991),
            .ce(),
            .sr(N__49115));
    defparam \phase_controller_inst1.test22_LC_12_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.test22_LC_12_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.test22_LC_12_6_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \phase_controller_inst1.test22_LC_12_6_4  (
            .in0(N__31027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30988),
            .lcout(test22_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49991),
            .ce(),
            .sr(N__49115));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_12_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_12_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_12_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_12_7_0  (
            .in0(N__50493),
            .in1(N__40249),
            .in2(_gnd_net_),
            .in3(N__43369),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49983),
            .ce(N__49465),
            .sr(N__49123));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_12_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_12_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_12_8_1  (
            .in0(N__31247),
            .in1(N__31178),
            .in2(N__31256),
            .in3(N__31241),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_12_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_12_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_12_8_6  (
            .in0(N__31305),
            .in1(N__34777),
            .in2(_gnd_net_),
            .in3(N__32189),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(N__32725),
            .sr(N__49130));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_12_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_12_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_12_9_0  (
            .in0(N__35275),
            .in1(N__35189),
            .in2(N__35526),
            .in3(N__34512),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_12_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_12_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_12_9_1  (
            .in0(N__34706),
            .in1(N__34565),
            .in2(N__34644),
            .in3(N__34766),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_12_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_12_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_12_9_2  (
            .in0(N__34100),
            .in1(N__34029),
            .in2(N__34173),
            .in3(N__34229),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_6  (
            .in0(N__31217),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31189),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_12_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_12_9_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_12_9_7  (
            .in0(N__34830),
            .in1(N__34998),
            .in2(N__34934),
            .in3(N__33960),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__31171),
            .in2(N__31136),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_12_10_1  (
            .in0(N__32704),
            .in1(N__31123),
            .in2(_gnd_net_),
            .in3(N__31109),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49958),
            .ce(),
            .sr(N__49142));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_12_10_2  (
            .in0(N__32722),
            .in1(N__31106),
            .in2(N__31099),
            .in3(N__31079),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49958),
            .ce(),
            .sr(N__49142));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_12_10_3  (
            .in0(N__32705),
            .in1(N__31474),
            .in2(_gnd_net_),
            .in3(N__31460),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49958),
            .ce(),
            .sr(N__49142));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_12_10_4  (
            .in0(N__32723),
            .in1(N__31453),
            .in2(_gnd_net_),
            .in3(N__31439),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49958),
            .ce(),
            .sr(N__49142));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_12_10_5  (
            .in0(N__32706),
            .in1(N__31432),
            .in2(_gnd_net_),
            .in3(N__31418),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49958),
            .ce(),
            .sr(N__49142));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_12_10_6  (
            .in0(N__32724),
            .in1(N__31411),
            .in2(_gnd_net_),
            .in3(N__31397),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49958),
            .ce(),
            .sr(N__49142));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_10_7  (
            .in0(N__32707),
            .in1(N__31390),
            .in2(_gnd_net_),
            .in3(N__31376),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49958),
            .ce(),
            .sr(N__49142));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_11_0  (
            .in0(N__32715),
            .in1(N__31369),
            .in2(_gnd_net_),
            .in3(N__31355),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49149));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_12_11_1  (
            .in0(N__32708),
            .in1(N__31348),
            .in2(_gnd_net_),
            .in3(N__31334),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49149));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_12_11_2  (
            .in0(N__32712),
            .in1(N__31327),
            .in2(_gnd_net_),
            .in3(N__31313),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49149));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_12_11_3  (
            .in0(N__32709),
            .in1(N__31663),
            .in2(_gnd_net_),
            .in3(N__31649),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49149));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_12_11_4  (
            .in0(N__32713),
            .in1(N__31642),
            .in2(_gnd_net_),
            .in3(N__31628),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49149));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_12_11_5  (
            .in0(N__32710),
            .in1(N__31621),
            .in2(_gnd_net_),
            .in3(N__31607),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49149));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_12_11_6  (
            .in0(N__32714),
            .in1(N__31600),
            .in2(_gnd_net_),
            .in3(N__31586),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49149));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_12_11_7  (
            .in0(N__32711),
            .in1(N__31573),
            .in2(_gnd_net_),
            .in3(N__31559),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49949),
            .ce(),
            .sr(N__49149));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_12_12_0  (
            .in0(N__32689),
            .in1(N__31554),
            .in2(_gnd_net_),
            .in3(N__31538),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_12_12_1  (
            .in0(N__32672),
            .in1(N__31525),
            .in2(_gnd_net_),
            .in3(N__31511),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_12_12_2  (
            .in0(N__32690),
            .in1(N__31495),
            .in2(_gnd_net_),
            .in3(N__31481),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_12_12_3  (
            .in0(N__32673),
            .in1(N__31896),
            .in2(_gnd_net_),
            .in3(N__31874),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_12_12_4  (
            .in0(N__32691),
            .in1(N__31866),
            .in2(_gnd_net_),
            .in3(N__31847),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_12_12_5  (
            .in0(N__32674),
            .in1(N__31837),
            .in2(_gnd_net_),
            .in3(N__31823),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_12_12_6  (
            .in0(N__32692),
            .in1(N__31806),
            .in2(_gnd_net_),
            .in3(N__31790),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_12_12_7  (
            .in0(N__32675),
            .in1(N__31779),
            .in2(_gnd_net_),
            .in3(N__31763),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49155));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_12_13_0  (
            .in0(N__32665),
            .in1(N__31753),
            .in2(_gnd_net_),
            .in3(N__31739),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49161));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_12_13_1  (
            .in0(N__32669),
            .in1(N__31731),
            .in2(_gnd_net_),
            .in3(N__31715),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49161));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_12_13_2  (
            .in0(N__32666),
            .in1(N__31710),
            .in2(_gnd_net_),
            .in3(N__31694),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49161));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_12_13_3  (
            .in0(N__32670),
            .in1(N__31686),
            .in2(_gnd_net_),
            .in3(N__31670),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49161));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_12_13_4  (
            .in0(N__32667),
            .in1(N__32790),
            .in2(_gnd_net_),
            .in3(N__32774),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49161));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_12_13_5  (
            .in0(N__32671),
            .in1(N__32760),
            .in2(_gnd_net_),
            .in3(N__32741),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49161));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_12_13_6  (
            .in0(N__32668),
            .in1(N__32472),
            .in2(_gnd_net_),
            .in3(N__32477),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49161));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_12_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_12_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_12_14_0  (
            .in0(N__32448),
            .in1(N__34566),
            .in2(_gnd_net_),
            .in3(N__32413),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_12_14_4  (
            .in0(N__34166),
            .in1(N__32001),
            .in2(_gnd_net_),
            .in3(N__32412),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_12_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_12_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_12_16_0 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_inst1.state_3_LC_12_16_0  (
            .in0(N__31975),
            .in1(N__35678),
            .in2(N__35887),
            .in3(N__31964),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49919),
            .ce(),
            .sr(N__49176));
    defparam \phase_controller_inst2.stoper_hc.running_LC_12_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_12_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_12_16_1 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_12_16_1  (
            .in0(N__31913),
            .in1(N__36682),
            .in2(N__31958),
            .in3(N__38391),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49919),
            .ce(),
            .sr(N__49176));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_16_2 .LUT_INIT=16'b0100111001001110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_12_16_2  (
            .in0(N__35704),
            .in1(N__36128),
            .in2(N__36164),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49919),
            .ce(),
            .sr(N__49176));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_12_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_12_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__32948),
            .in2(N__32942),
            .in3(N__32934),
            .lcout(\current_shift_inst.control_input_1 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_17_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__35582),
            .in2(_gnd_net_),
            .in3(N__32897),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_17_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__35576),
            .in2(_gnd_net_),
            .in3(N__32882),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__35570),
            .in2(_gnd_net_),
            .in3(N__32870),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_17_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__35564),
            .in2(_gnd_net_),
            .in3(N__32858),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_17_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__35765),
            .in2(_gnd_net_),
            .in3(N__32843),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_17_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__35759),
            .in2(_gnd_net_),
            .in3(N__32831),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_17_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__35711),
            .in2(_gnd_net_),
            .in3(N__32816),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_18_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__32813),
            .in2(_gnd_net_),
            .in3(N__32795),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_18_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33065),
            .in3(N__33047),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_18_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__35594),
            .in2(_gnd_net_),
            .in3(N__33032),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_18_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__38867),
            .in2(_gnd_net_),
            .in3(N__33020),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_18_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__38894),
            .in2(_gnd_net_),
            .in3(N__33008),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_18_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__39059),
            .in2(_gnd_net_),
            .in3(N__32993),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_12 ),
            .carryout(\current_shift_inst.control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_12_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_12_18_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__39032),
            .in2(_gnd_net_),
            .in3(N__32981),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_13 ),
            .carryout(\current_shift_inst.control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_12_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_12_18_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(N__39008),
            .in2(_gnd_net_),
            .in3(N__32966),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_14 ),
            .carryout(\current_shift_inst.control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_12_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_12_19_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__35588),
            .in2(_gnd_net_),
            .in3(N__32951),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\current_shift_inst.control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_12_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_12_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__35747),
            .in2(_gnd_net_),
            .in3(N__33164),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_16 ),
            .carryout(\current_shift_inst.control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_12_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_12_19_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(N__35753),
            .in2(_gnd_net_),
            .in3(N__33149),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_17 ),
            .carryout(\current_shift_inst.control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_12_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_12_19_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__37232),
            .in2(_gnd_net_),
            .in3(N__33137),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_18 ),
            .carryout(\current_shift_inst.control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_12_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_12_19_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__35741),
            .in2(_gnd_net_),
            .in3(N__33125),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_19 ),
            .carryout(\current_shift_inst.control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_12_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_12_19_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(N__35735),
            .in2(_gnd_net_),
            .in3(N__33110),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_20 ),
            .carryout(\current_shift_inst.control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_12_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_12_19_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__35729),
            .in2(_gnd_net_),
            .in3(N__33098),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_21 ),
            .carryout(\current_shift_inst.control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_12_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_12_19_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__39152),
            .in2(_gnd_net_),
            .in3(N__33083),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_22 ),
            .carryout(\current_shift_inst.control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_12_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_12_20_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__38843),
            .in2(_gnd_net_),
            .in3(N__33068),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\current_shift_inst.control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_12_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_12_20_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__36008),
            .in2(_gnd_net_),
            .in3(N__33305),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_24 ),
            .carryout(\current_shift_inst.control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_12_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_12_20_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__35717),
            .in2(_gnd_net_),
            .in3(N__33290),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_25 ),
            .carryout(\current_shift_inst.control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_12_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_12_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__35723),
            .in2(_gnd_net_),
            .in3(N__33278),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_26 ),
            .carryout(\current_shift_inst.control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_12_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_12_20_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__37145),
            .in2(_gnd_net_),
            .in3(N__33266),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_27 ),
            .carryout(\current_shift_inst.control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_12_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_12_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__36002),
            .in2(_gnd_net_),
            .in3(N__33251),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_28 ),
            .carryout(\current_shift_inst.control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_12_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_12_20_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__41873),
            .in2(_gnd_net_),
            .in3(N__33248),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_12_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_12_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33241),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1  (
            .in0(N__49268),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_13_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_13_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_13_4_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \phase_controller_inst1.state_1_LC_13_4_0  (
            .in0(N__33386),
            .in1(N__33212),
            .in2(_gnd_net_),
            .in3(N__35798),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50028),
            .ce(),
            .sr(N__49100));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_4_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_4_1  (
            .in0(N__39450),
            .in1(N__39476),
            .in2(N__37345),
            .in3(N__49429),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50028),
            .ce(),
            .sr(N__49100));
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_4_4 .LUT_INIT=16'b1011111100001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_13_4_4  (
            .in0(N__39505),
            .in1(N__39451),
            .in2(N__39549),
            .in3(N__39271),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50028),
            .ce(),
            .sr(N__49100));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39251),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50028),
            .ce(),
            .sr(N__49100));
    defparam \phase_controller_inst1.start_timer_hc_LC_13_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_4_7 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_13_4_7  (
            .in0(N__33395),
            .in1(N__33385),
            .in2(N__39257),
            .in3(N__33370),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50028),
            .ce(),
            .sr(N__49100));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_13_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_13_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_13_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_13_5_1  (
            .in0(N__39228),
            .in1(N__42671),
            .in2(_gnd_net_),
            .in3(N__50496),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50015),
            .ce(N__49543),
            .sr(N__49105));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_13_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_13_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_13_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_13_5_5  (
            .in0(N__44387),
            .in1(N__44340),
            .in2(_gnd_net_),
            .in3(N__50495),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50015),
            .ce(N__49543),
            .sr(N__49105));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_5_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_13_5_6  (
            .in0(N__50494),
            .in1(N__37937),
            .in2(_gnd_net_),
            .in3(N__42389),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50015),
            .ce(N__49543),
            .sr(N__49105));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_13_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_13_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_13_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_13_5_7  (
            .in0(N__42524),
            .in1(N__37912),
            .in2(_gnd_net_),
            .in3(N__50497),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50015),
            .ce(N__49543),
            .sr(N__49105));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_13_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_13_6_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_13_6_1  (
            .in0(N__36316),
            .in1(N__37799),
            .in2(N__36344),
            .in3(N__37826),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_13_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_13_6_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_13_6_4  (
            .in0(N__50481),
            .in1(N__44341),
            .in2(_gnd_net_),
            .in3(N__44386),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_13_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_13_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_13_6_5  (
            .in0(N__42573),
            .in1(N__37948),
            .in2(_gnd_net_),
            .in3(N__50482),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(elapsed_time_ns_1_RNIH33T9_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_13_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_13_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_13_6_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_13_6_6  (
            .in0(N__50483),
            .in1(_gnd_net_),
            .in2(N__33401),
            .in3(N__42574),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50005),
            .ce(N__49500),
            .sr(N__49110));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_6_7  (
            .in0(N__44298),
            .in1(N__44272),
            .in2(_gnd_net_),
            .in3(N__50480),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_7_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_7_0  (
            .in0(N__36383),
            .in1(N__37856),
            .in2(N__37613),
            .in3(N__36371),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_13_7_1  (
            .in0(N__50485),
            .in1(N__40276),
            .in2(_gnd_net_),
            .in3(N__43425),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_13_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_13_7_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_13_7_2  (
            .in0(N__43426),
            .in1(_gnd_net_),
            .in2(N__33398),
            .in3(N__50486),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49994),
            .ce(N__49577),
            .sr(N__49116));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_13_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_13_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_13_8_1  (
            .in0(N__36459),
            .in1(N__43555),
            .in2(_gnd_net_),
            .in3(N__50522),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49984),
            .ce(N__49549),
            .sr(N__49124));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_13_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_13_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_13_8_7  (
            .in0(N__43985),
            .in1(N__37872),
            .in2(_gnd_net_),
            .in3(N__50523),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49984),
            .ce(N__49549),
            .sr(N__49124));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_13_9_1  (
            .in0(N__37936),
            .in1(N__42388),
            .in2(_gnd_net_),
            .in3(N__50526),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__35663),
            .in2(_gnd_net_),
            .in3(N__35888),
            .lcout(\phase_controller_inst1.test_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__33790),
            .in2(N__33938),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49968),
            .ce(N__35105),
            .sr(N__49137));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__33712),
            .in2(N__33869),
            .in3(N__33794),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49968),
            .ce(N__35105),
            .sr(N__49137));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__33791),
            .in2(N__33644),
            .in3(N__33719),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49968),
            .ce(N__35105),
            .sr(N__49137));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__33568),
            .in2(N__33716),
            .in3(N__33647),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49968),
            .ce(N__35105),
            .sr(N__49137));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__33643),
            .in2(N__33502),
            .in3(N__33575),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49968),
            .ce(N__35105),
            .sr(N__49137));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__33424),
            .in2(N__33572),
            .in3(N__33506),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49968),
            .ce(N__35105),
            .sr(N__49137));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__34429),
            .in2(N__33503),
            .in3(N__33431),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49968),
            .ce(N__35105),
            .sr(N__49137));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__34348),
            .in2(N__33428),
            .in3(N__34439),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49968),
            .ce(N__35105),
            .sr(N__49137));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__34267),
            .in2(N__34436),
            .in3(N__34355),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49961),
            .ce(N__35104),
            .sr(N__49143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__34198),
            .in2(N__34352),
            .in3(N__34274),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49961),
            .ce(N__35104),
            .sr(N__49143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__34129),
            .in2(N__34271),
            .in3(N__34205),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49961),
            .ce(N__35104),
            .sr(N__49143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__34069),
            .in2(N__34202),
            .in3(N__34136),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49961),
            .ce(N__35104),
            .sr(N__49143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__33997),
            .in2(N__34133),
            .in3(N__34076),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49961),
            .ce(N__35104),
            .sr(N__49143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__35035),
            .in2(N__34073),
            .in3(N__34004),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49961),
            .ce(N__35104),
            .sr(N__49143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__34972),
            .in2(N__34001),
            .in3(N__33941),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49961),
            .ce(N__35104),
            .sr(N__49143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__35036),
            .in2(N__34891),
            .in3(N__34982),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49961),
            .ce(N__35104),
            .sr(N__49143));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__34807),
            .in2(N__34979),
            .in3(N__34895),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49952),
            .ce(N__35100),
            .sr(N__49150));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__34741),
            .in2(N__34892),
            .in3(N__34814),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49952),
            .ce(N__35100),
            .sr(N__49150));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__34669),
            .in2(N__34811),
            .in3(N__34748),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49952),
            .ce(N__35100),
            .sr(N__49150));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__34597),
            .in2(N__34745),
            .in3(N__34676),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49952),
            .ce(N__35100),
            .sr(N__49150));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__34534),
            .in2(N__34673),
            .in3(N__34601),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49952),
            .ce(N__35100),
            .sr(N__49150));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__34598),
            .in2(N__35557),
            .in3(N__34538),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49952),
            .ce(N__35100),
            .sr(N__49150));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__34535),
            .in2(N__35480),
            .in3(N__34472),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49952),
            .ce(N__35100),
            .sr(N__49150));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__35398),
            .in2(N__35558),
            .in3(N__35483),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49952),
            .ce(N__35100),
            .sr(N__49150));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__35299),
            .in2(N__35479),
            .in3(N__35402),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49945),
            .ce(N__35086),
            .sr(N__49156));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__35399),
            .in2(N__35218),
            .in3(N__35324),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49945),
            .ce(N__35086),
            .sr(N__49156));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__35321),
            .in2(N__35303),
            .in3(N__35240),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49945),
            .ce(N__35086),
            .sr(N__49156));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__35237),
            .in2(N__35219),
            .in3(N__35156),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49945),
            .ce(N__35086),
            .sr(N__49156));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35153),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(N__35086),
            .sr(N__49156));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(N__35705),
            .in2(_gnd_net_),
            .in3(N__36156),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_163_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_15_5 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_13_15_5  (
            .in0(N__36157),
            .in1(N__35700),
            .in2(_gnd_net_),
            .in3(N__36124),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_164_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_16_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_16_0  (
            .in0(N__38594),
            .in1(N__37025),
            .in2(_gnd_net_),
            .in3(N__41837),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35699),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.test_LC_13_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.test_LC_13_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.test_LC_13_17_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \phase_controller_inst1.test_LC_13_17_5  (
            .in0(N__35671),
            .in1(N__35605),
            .in2(_gnd_net_),
            .in3(N__35874),
            .lcout(test_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49921),
            .ce(),
            .sr(N__49177));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_13_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_13_18_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_13_18_0  (
            .in0(N__38549),
            .in1(N__36986),
            .in2(_gnd_net_),
            .in3(N__41810),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_18_1 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_18_1  (
            .in0(N__41811),
            .in1(_gnd_net_),
            .in2(N__38735),
            .in3(N__37115),
            .lcout(\current_shift_inst.control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_13_18_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_13_18_2  (
            .in0(N__36938),
            .in1(N__38498),
            .in2(_gnd_net_),
            .in3(N__41804),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_13_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_13_18_3 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_13_18_3  (
            .in0(N__41805),
            .in1(_gnd_net_),
            .in2(N__38480),
            .in3(N__36926),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_13_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_13_18_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_13_18_4  (
            .in0(N__38462),
            .in1(N__36911),
            .in2(_gnd_net_),
            .in3(N__41806),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_13_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_13_18_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_13_18_5  (
            .in0(N__41807),
            .in1(N__38447),
            .in2(_gnd_net_),
            .in3(N__37064),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_18_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_18_6  (
            .in0(N__37049),
            .in1(N__38624),
            .in2(_gnd_net_),
            .in3(N__41808),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_18_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_18_7  (
            .in0(N__41809),
            .in1(N__38609),
            .in2(_gnd_net_),
            .in3(N__37037),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_19_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_19_0  (
            .in0(N__41865),
            .in1(N__37094),
            .in2(_gnd_net_),
            .in3(N__38699),
            .lcout(\current_shift_inst.control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_19_1 .LUT_INIT=16'b0101010100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_19_1  (
            .in0(N__37106),
            .in1(_gnd_net_),
            .in2(N__38717),
            .in3(N__41864),
            .lcout(\current_shift_inst.control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_19_2  (
            .in0(N__41866),
            .in1(_gnd_net_),
            .in2(N__38669),
            .in3(N__37076),
            .lcout(\current_shift_inst.control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_19_3  (
            .in0(N__38651),
            .in1(N__37199),
            .in2(_gnd_net_),
            .in3(N__41867),
            .lcout(\current_shift_inst.control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_19_4  (
            .in0(N__41868),
            .in1(N__37190),
            .in2(_gnd_net_),
            .in3(N__38636),
            .lcout(\current_shift_inst.control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_19_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_19_5  (
            .in0(N__38786),
            .in1(N__37157),
            .in2(_gnd_net_),
            .in3(N__41871),
            .lcout(\current_shift_inst.control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_19_6  (
            .in0(N__41870),
            .in1(N__38804),
            .in2(_gnd_net_),
            .in3(N__37166),
            .lcout(\current_shift_inst.control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_19_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_19_7  (
            .in0(N__38822),
            .in1(N__37175),
            .in2(_gnd_net_),
            .in3(N__41869),
            .lcout(\current_shift_inst.control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41872),
            .lcout(\current_shift_inst.control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35957),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35933),
            .ce(),
            .sr(N__49198));
    defparam \delay_measurement_inst.start_timer_tr_LC_13_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_13_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_13_21_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_13_21_5  (
            .in0(N__35958),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35933),
            .ce(),
            .sr(N__49198));
    defparam \current_shift_inst.stop_timer_s1_LC_13_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_13_22_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_22_0  (
            .in0(N__37463),
            .in1(N__35889),
            .in2(N__37421),
            .in3(N__35911),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49203));
    defparam \phase_controller_inst1.S1_LC_13_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_22_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.S1_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__35890),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49203));
    defparam \current_shift_inst.start_timer_s1_LC_13_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_13_23_4 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_23_4  (
            .in0(N__35910),
            .in1(N__37461),
            .in2(_gnd_net_),
            .in3(N__35894),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49899),
            .ce(),
            .sr(N__49206));
    defparam \current_shift_inst.timer_s1.running_LC_13_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_23_7 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_23_7  (
            .in0(N__37462),
            .in1(N__37416),
            .in2(_gnd_net_),
            .in3(N__37442),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49899),
            .ce(),
            .sr(N__49206));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__37420),
            .in2(_gnd_net_),
            .in3(N__37439),
            .lcout(\current_shift_inst.timer_s1.N_161_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_28_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_28_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35824),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49894),
            .ce(),
            .sr(N__49232));
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_3_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_3_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_14_3_0  (
            .in0(N__36109),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(),
            .sr(N__49091));
    defparam \delay_measurement_inst.start_timer_hc_LC_14_3_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_14_3_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_14_3_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_14_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36108),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36092),
            .ce(),
            .sr(N__49091));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_14_4_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_14_4_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_14_4_0  (
            .in0(N__37335),
            .in1(N__37370),
            .in2(N__36083),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_14_4_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_14_4_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_14_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(N__37382),
            .in2(N__36074),
            .in3(N__37319),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_14_4_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_14_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_14_4_2  (
            .in0(_gnd_net_),
            .in1(N__36065),
            .in2(N__36059),
            .in3(N__37300),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_14_4_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_14_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_14_4_3  (
            .in0(_gnd_net_),
            .in1(N__37376),
            .in2(N__36050),
            .in3(N__37582),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_14_4_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_14_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_14_4_4  (
            .in0(_gnd_net_),
            .in1(N__36041),
            .in2(N__36032),
            .in3(N__37567),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_14_4_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_14_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_14_4_5  (
            .in0(_gnd_net_),
            .in1(N__36014),
            .in2(N__36023),
            .in3(N__37552),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_14_4_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_14_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_14_4_6  (
            .in0(_gnd_net_),
            .in1(N__36245),
            .in2(N__37391),
            .in3(N__37537),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_14_4_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_14_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_14_4_7  (
            .in0(_gnd_net_),
            .in1(N__36239),
            .in2(N__36233),
            .in3(N__37522),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_14_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_14_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(N__41108),
            .in2(N__36224),
            .in3(N__37507),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_14_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_14_5_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_14_5_1  (
            .in0(N__37492),
            .in1(N__41075),
            .in2(N__36215),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_14_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_14_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__41039),
            .in2(N__36206),
            .in3(N__37477),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_14_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_14_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(N__42683),
            .in2(N__36197),
            .in3(N__37723),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_14_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_14_5_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_14_5_4  (
            .in0(N__37708),
            .in1(N__39794),
            .in2(N__36185),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_14_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_14_5_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_14_5_5  (
            .in0(N__37693),
            .in1(N__40820),
            .in2(N__36176),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_14_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_14_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__36470),
            .in2(N__36269),
            .in3(N__37678),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_14_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_14_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__40913),
            .in2(N__40985),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_14_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_14_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__36350),
            .in2(N__36281),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_14_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_14_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__36356),
            .in2(N__36260),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_14_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_14_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__39680),
            .in2(N__39635),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_14_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_14_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__36251),
            .in2(N__36305),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_14_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_14_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__36389),
            .in2(N__36407),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_14_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_14_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__39356),
            .in2(N__39413),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_14_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_14_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(N__39806),
            .in2(N__39590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36410),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_14_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_14_7_0 .LUT_INIT=16'b0111010100010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_14_7_0  (
            .in0(N__37746),
            .in1(N__37764),
            .in2(N__37364),
            .in3(N__36398),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_14_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_14_7_1 .LUT_INIT=16'b1000101011101111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_14_7_1  (
            .in0(N__36397),
            .in1(N__37363),
            .in2(N__37769),
            .in3(N__37747),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_14_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_14_7_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_14_7_2  (
            .in0(N__36382),
            .in1(N__37851),
            .in2(N__37612),
            .in3(N__36370),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_14_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_14_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_14_7_4  (
            .in0(N__37876),
            .in1(N__43984),
            .in2(_gnd_net_),
            .in3(N__50500),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_14_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_14_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_14_7_5  (
            .in0(N__50499),
            .in1(N__42513),
            .in2(_gnd_net_),
            .in3(N__37911),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_14_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_14_7_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_14_7_6  (
            .in0(N__36296),
            .in1(N__37633),
            .in2(N__37658),
            .in3(N__36487),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_7_7 .LUT_INIT=16'b0010101100001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_7_7  (
            .in0(N__36343),
            .in1(N__37821),
            .in2(N__37798),
            .in3(N__36320),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_8_0 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_8_0  (
            .in0(N__36292),
            .in1(N__37653),
            .in2(N__36488),
            .in3(N__37632),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_14_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_14_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_14_8_1  (
            .in0(N__43554),
            .in1(N__36461),
            .in2(_gnd_net_),
            .in3(N__50394),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_14_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_14_8_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_14_8_2  (
            .in0(N__43489),
            .in1(_gnd_net_),
            .in2(N__50498),
            .in3(N__36433),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(elapsed_time_ns_1_RNI68CN9_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_14_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_14_8_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__43490),
            .in2(N__36491),
            .in3(N__50396),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49995),
            .ce(N__49548),
            .sr(N__49117));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_8_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_8_5  (
            .in0(N__42867),
            .in1(N__50390),
            .in2(_gnd_net_),
            .in3(N__37888),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(elapsed_time_ns_1_RNI24CN9_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_14_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_14_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_14_8_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_14_8_6  (
            .in0(N__50395),
            .in1(_gnd_net_),
            .in2(N__36473),
            .in3(N__42868),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49995),
            .ce(N__49548),
            .sr(N__49117));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_9_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_14_9_0  (
            .in0(N__36614),
            .in1(N__36637),
            .in2(N__36422),
            .in3(N__36443),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_14_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_14_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_14_9_1  (
            .in0(N__36442),
            .in1(N__36613),
            .in2(N__36641),
            .in3(N__36418),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_14_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_14_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_14_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_14_9_2  (
            .in0(N__36460),
            .in1(N__43559),
            .in2(_gnd_net_),
            .in3(N__50518),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49985),
            .ce(N__45112),
            .sr(N__49125));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_14_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_14_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_14_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_14_9_3  (
            .in0(N__50516),
            .in1(N__43488),
            .in2(_gnd_net_),
            .in3(N__36434),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49985),
            .ce(N__45112),
            .sr(N__49125));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_14_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_14_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_14_9_4  (
            .in0(N__39233),
            .in1(N__42670),
            .in2(_gnd_net_),
            .in3(N__50519),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49985),
            .ce(N__45112),
            .sr(N__49125));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_14_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_14_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_14_9_5  (
            .in0(N__50517),
            .in1(N__39299),
            .in2(_gnd_net_),
            .in3(N__42635),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49985),
            .ce(N__45112),
            .sr(N__49125));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__36548),
            .in2(N__38162),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_14_10_1  (
            .in0(N__36874),
            .in1(N__38120),
            .in2(_gnd_net_),
            .in3(N__36530),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49975),
            .ce(),
            .sr(N__49131));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_14_10_2  (
            .in0(N__36878),
            .in1(N__38089),
            .in2(N__36527),
            .in3(N__36506),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49975),
            .ce(),
            .sr(N__49131));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_14_10_3  (
            .in0(N__36875),
            .in1(N__38069),
            .in2(_gnd_net_),
            .in3(N__36503),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49975),
            .ce(),
            .sr(N__49131));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_14_10_4  (
            .in0(N__36879),
            .in1(N__38036),
            .in2(_gnd_net_),
            .in3(N__36500),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49975),
            .ce(),
            .sr(N__49131));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_14_10_5  (
            .in0(N__36876),
            .in1(N__38012),
            .in2(_gnd_net_),
            .in3(N__36497),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49975),
            .ce(),
            .sr(N__49131));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_14_10_6  (
            .in0(N__36880),
            .in1(N__37981),
            .in2(_gnd_net_),
            .in3(N__36494),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49975),
            .ce(),
            .sr(N__49131));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_14_10_7  (
            .in0(N__36877),
            .in1(N__38345),
            .in2(_gnd_net_),
            .in3(N__36575),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49975),
            .ce(),
            .sr(N__49131));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_14_11_0  (
            .in0(N__36866),
            .in1(N__38324),
            .in2(_gnd_net_),
            .in3(N__36572),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49969),
            .ce(),
            .sr(N__49138));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_14_11_1  (
            .in0(N__36831),
            .in1(N__38303),
            .in2(_gnd_net_),
            .in3(N__36569),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49969),
            .ce(),
            .sr(N__49138));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_14_11_2  (
            .in0(N__36863),
            .in1(N__38282),
            .in2(_gnd_net_),
            .in3(N__36566),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49969),
            .ce(),
            .sr(N__49138));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_14_11_3  (
            .in0(N__36832),
            .in1(N__38261),
            .in2(_gnd_net_),
            .in3(N__36563),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49969),
            .ce(),
            .sr(N__49138));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_14_11_4  (
            .in0(N__36864),
            .in1(N__38240),
            .in2(_gnd_net_),
            .in3(N__36560),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49969),
            .ce(),
            .sr(N__49138));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_14_11_5  (
            .in0(N__36833),
            .in1(N__38219),
            .in2(_gnd_net_),
            .in3(N__36557),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49969),
            .ce(),
            .sr(N__49138));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_14_11_6  (
            .in0(N__36865),
            .in1(N__38189),
            .in2(_gnd_net_),
            .in3(N__36554),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49969),
            .ce(),
            .sr(N__49138));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_14_11_7  (
            .in0(N__36834),
            .in1(N__39766),
            .in2(_gnd_net_),
            .in3(N__36551),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49969),
            .ce(),
            .sr(N__49138));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_14_12_0  (
            .in0(N__36851),
            .in1(N__39742),
            .in2(_gnd_net_),
            .in3(N__36644),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49144));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_14_12_1  (
            .in0(N__36855),
            .in1(N__36631),
            .in2(_gnd_net_),
            .in3(N__36617),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49144));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_14_12_2  (
            .in0(N__36852),
            .in1(N__36612),
            .in2(_gnd_net_),
            .in3(N__36596),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49144));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_14_12_3  (
            .in0(N__36856),
            .in1(N__40303),
            .in2(_gnd_net_),
            .in3(N__36593),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49144));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_14_12_4  (
            .in0(N__36853),
            .in1(N__40327),
            .in2(_gnd_net_),
            .in3(N__36590),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49144));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_14_12_5  (
            .in0(N__36857),
            .in1(N__40164),
            .in2(_gnd_net_),
            .in3(N__36587),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49144));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_14_12_6  (
            .in0(N__36854),
            .in1(N__40147),
            .in2(_gnd_net_),
            .in3(N__36584),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49144));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_14_12_7  (
            .in0(N__36858),
            .in1(N__44436),
            .in2(_gnd_net_),
            .in3(N__36581),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49962),
            .ce(),
            .sr(N__49144));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_14_13_0  (
            .in0(N__36859),
            .in1(N__44410),
            .in2(_gnd_net_),
            .in3(N__36578),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49953),
            .ce(),
            .sr(N__49151));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_14_13_1  (
            .in0(N__36867),
            .in1(N__40027),
            .in2(_gnd_net_),
            .in3(N__36899),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49953),
            .ce(),
            .sr(N__49151));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_14_13_2  (
            .in0(N__36860),
            .in1(N__40063),
            .in2(_gnd_net_),
            .in3(N__36896),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49953),
            .ce(),
            .sr(N__49151));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_14_13_3  (
            .in0(N__36868),
            .in1(N__39937),
            .in2(_gnd_net_),
            .in3(N__36893),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49953),
            .ce(),
            .sr(N__49151));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_14_13_4  (
            .in0(N__36861),
            .in1(N__39913),
            .in2(_gnd_net_),
            .in3(N__36890),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49953),
            .ce(),
            .sr(N__49151));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_14_13_5  (
            .in0(N__36869),
            .in1(N__44191),
            .in2(_gnd_net_),
            .in3(N__36887),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49953),
            .ce(),
            .sr(N__49151));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_14_13_6  (
            .in0(N__36862),
            .in1(N__44167),
            .in2(_gnd_net_),
            .in3(N__36884),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49953),
            .ce(),
            .sr(N__49151));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_13_7 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_14_13_7  (
            .in0(N__36870),
            .in1(N__36728),
            .in2(N__36701),
            .in3(N__38157),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49953),
            .ce(),
            .sr(N__49151));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_14_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_14_14_4  (
            .in0(N__46375),
            .in1(N__45832),
            .in2(N__46880),
            .in3(N__40582),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__47758),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49946),
            .ce(N__47792),
            .sr(N__49157));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_14_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_14_14_6  (
            .in0(N__46376),
            .in1(N__45833),
            .in2(N__46879),
            .in3(N__40583),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_7  (
            .in0(N__45831),
            .in1(N__46377),
            .in2(N__46930),
            .in3(N__40613),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__44627),
            .in2(N__45653),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_15_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_15_1  (
            .in0(N__45023),
            .in1(N__40473),
            .in2(N__40505),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__46252),
            .in2(N__36968),
            .in3(N__45024),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__36959),
            .in2(N__46439),
            .in3(N__36941),
            .lcout(\current_shift_inst.un38_control_input_0_s0_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__46256),
            .in2(N__41315),
            .in3(N__36929),
            .lcout(\current_shift_inst.un38_control_input_0_s0_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__44525),
            .in2(N__46440),
            .in3(N__36914),
            .lcout(\current_shift_inst.un38_control_input_0_s0_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__46260),
            .in2(N__38948),
            .in3(N__36902),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__37133),
            .in2(N__46441),
            .in3(N__37052),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__46280),
            .in2(N__46673),
            .in3(N__37040),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__40559),
            .in2(N__46446),
            .in3(N__37028),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__46284),
            .in2(N__46058),
            .in3(N__37019),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__38753),
            .in2(N__46447),
            .in3(N__37004),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__46288),
            .in2(N__41651),
            .in3(N__36989),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__38747),
            .in2(N__46448),
            .in3(N__36977),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__46292),
            .in2(N__38933),
            .in3(N__36974),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__45179),
            .in2(N__46449),
            .in3(N__36971),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__46450),
            .in2(N__41378),
            .in3(N__37124),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__37217),
            .in2(N__46593),
            .in3(N__37121),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__46454),
            .in2(N__37262),
            .in3(N__37118),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__38999),
            .in2(N__46594),
            .in3(N__37109),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__46458),
            .in2(N__37286),
            .in3(N__37097),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__38993),
            .in2(N__46595),
            .in3(N__37082),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__46462),
            .in2(N__37274),
            .in3(N__37079),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__37250),
            .in2(N__46596),
            .in3(N__37067),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__37223),
            .in2(N__46597),
            .in3(N__37193),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__46469),
            .in2(N__39194),
            .in3(N__37184),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__38954),
            .in2(N__46598),
            .in3(N__37181),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__46473),
            .in2(N__39176),
            .in3(N__37178),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__37208),
            .in2(N__46599),
            .in3(N__37169),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__46477),
            .in2(N__39143),
            .in3(N__37160),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__39332),
            .in2(N__46600),
            .in3(N__37151),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_18_7 .LUT_INIT=16'b1100010100110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_18_7  (
            .in0(N__38768),
            .in1(N__40541),
            .in2(N__41863),
            .in3(N__37148),
            .lcout(\current_shift_inst.control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_14_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_14_19_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_14_19_0  (
            .in0(N__45874),
            .in1(N__46561),
            .in2(N__47305),
            .in3(N__40708),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_19_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_19_1  (
            .in0(N__46564),
            .in1(N__45877),
            .in2(N__47474),
            .in3(N__45473),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_19_2  (
            .in0(N__45878),
            .in1(N__46562),
            .in2(N__42185),
            .in3(N__47383),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_3  (
            .in0(N__46560),
            .in1(N__45876),
            .in2(N__41924),
            .in3(N__47554),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4  (
            .in0(N__45879),
            .in1(N__46563),
            .in2(N__47345),
            .in3(N__45170),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_19_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_19_5  (
            .in0(N__38684),
            .in1(N__37241),
            .in2(_gnd_net_),
            .in3(N__41861),
            .lcout(\current_shift_inst.control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_19_6  (
            .in0(N__45880),
            .in1(N__46565),
            .in2(N__48059),
            .in3(N__42056),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_14_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_14_19_7 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_14_19_7  (
            .in0(N__46566),
            .in1(N__47599),
            .in2(N__45638),
            .in3(N__45875),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0  (
            .in0(N__45955),
            .in1(N__47876),
            .in2(N__46651),
            .in3(N__41720),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37440),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_23_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_23_4  (
            .in0(N__37460),
            .in1(N__37441),
            .in2(_gnd_net_),
            .in3(N__37415),
            .lcout(\current_shift_inst.timer_s1.N_162_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_15_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_15_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_15_4_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_15_4_0  (
            .in0(N__50477),
            .in1(N__40216),
            .in2(_gnd_net_),
            .in3(N__42455),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50042),
            .ce(N__49565),
            .sr(N__49092));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_15_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_15_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_15_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_15_4_1  (
            .in0(N__39567),
            .in1(N__43701),
            .in2(_gnd_net_),
            .in3(N__50479),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50042),
            .ce(N__49565),
            .sr(N__49092));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_15_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_15_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_15_4_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_15_4_2  (
            .in0(N__39288),
            .in1(_gnd_net_),
            .in2(N__50525),
            .in3(N__42631),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50042),
            .ce(N__49565),
            .sr(N__49092));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_15_4_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_15_4_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_15_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_15_4_3  (
            .in0(N__44480),
            .in1(N__44516),
            .in2(_gnd_net_),
            .in3(N__50478),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50042),
            .ce(N__49565),
            .sr(N__49092));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_15_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_15_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_15_4_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_15_4_4  (
            .in0(N__50473),
            .in1(N__39996),
            .in2(_gnd_net_),
            .in3(N__44063),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50042),
            .ce(N__49565),
            .sr(N__49092));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_15_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_15_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(N__39419),
            .in2(N__37349),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_5_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1  (
            .in0(N__49356),
            .in1(N__37318),
            .in2(_gnd_net_),
            .in3(N__37304),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__50036),
            .ce(),
            .sr(N__49095));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2  (
            .in0(N__49387),
            .in1(N__37301),
            .in2(N__39206),
            .in3(N__37289),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__50036),
            .ce(),
            .sr(N__49095));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3  (
            .in0(N__49357),
            .in1(N__37583),
            .in2(_gnd_net_),
            .in3(N__37571),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__50036),
            .ce(),
            .sr(N__49095));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4  (
            .in0(N__49388),
            .in1(N__37568),
            .in2(_gnd_net_),
            .in3(N__37556),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__50036),
            .ce(),
            .sr(N__49095));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5  (
            .in0(N__49358),
            .in1(N__37553),
            .in2(_gnd_net_),
            .in3(N__37541),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__50036),
            .ce(),
            .sr(N__49095));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6  (
            .in0(N__49389),
            .in1(N__37538),
            .in2(_gnd_net_),
            .in3(N__37526),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__50036),
            .ce(),
            .sr(N__49095));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7  (
            .in0(N__49359),
            .in1(N__37523),
            .in2(_gnd_net_),
            .in3(N__37511),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__50036),
            .ce(),
            .sr(N__49095));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0  (
            .in0(N__49525),
            .in1(N__37508),
            .in2(_gnd_net_),
            .in3(N__37496),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__50029),
            .ce(),
            .sr(N__49101));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1  (
            .in0(N__49433),
            .in1(N__37493),
            .in2(_gnd_net_),
            .in3(N__37481),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__50029),
            .ce(),
            .sr(N__49101));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2  (
            .in0(N__49522),
            .in1(N__37478),
            .in2(_gnd_net_),
            .in3(N__37466),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__50029),
            .ce(),
            .sr(N__49101));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3  (
            .in0(N__49434),
            .in1(N__37724),
            .in2(_gnd_net_),
            .in3(N__37712),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__50029),
            .ce(),
            .sr(N__49101));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4  (
            .in0(N__49523),
            .in1(N__37709),
            .in2(_gnd_net_),
            .in3(N__37697),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__50029),
            .ce(),
            .sr(N__49101));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5  (
            .in0(N__49435),
            .in1(N__37694),
            .in2(_gnd_net_),
            .in3(N__37682),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__50029),
            .ce(),
            .sr(N__49101));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6  (
            .in0(N__49524),
            .in1(N__37679),
            .in2(_gnd_net_),
            .in3(N__37667),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__50029),
            .ce(),
            .sr(N__49101));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7  (
            .in0(N__49436),
            .in1(N__40927),
            .in2(_gnd_net_),
            .in3(N__37664),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__50029),
            .ce(),
            .sr(N__49101));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0  (
            .in0(N__49526),
            .in1(N__40953),
            .in2(_gnd_net_),
            .in3(N__37661),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__50016),
            .ce(),
            .sr(N__49106));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1  (
            .in0(N__49461),
            .in1(N__37657),
            .in2(_gnd_net_),
            .in3(N__37637),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__50016),
            .ce(),
            .sr(N__49106));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2  (
            .in0(N__49527),
            .in1(N__37634),
            .in2(_gnd_net_),
            .in3(N__37616),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__50016),
            .ce(),
            .sr(N__49106));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3  (
            .in0(N__49462),
            .in1(N__37608),
            .in2(_gnd_net_),
            .in3(N__37586),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__50016),
            .ce(),
            .sr(N__49106));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4  (
            .in0(N__49528),
            .in1(N__37855),
            .in2(_gnd_net_),
            .in3(N__37835),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__50016),
            .ce(),
            .sr(N__49106));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5  (
            .in0(N__49463),
            .in1(N__39652),
            .in2(_gnd_net_),
            .in3(N__37832),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__50016),
            .ce(),
            .sr(N__49106));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6  (
            .in0(N__49529),
            .in1(N__39668),
            .in2(_gnd_net_),
            .in3(N__37829),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__50016),
            .ce(),
            .sr(N__49106));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7  (
            .in0(N__49464),
            .in1(N__37822),
            .in2(_gnd_net_),
            .in3(N__37802),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__50016),
            .ce(),
            .sr(N__49106));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0  (
            .in0(N__49469),
            .in1(N__37794),
            .in2(_gnd_net_),
            .in3(N__37772),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__50006),
            .ce(),
            .sr(N__49111));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1  (
            .in0(N__49578),
            .in1(N__37768),
            .in2(_gnd_net_),
            .in3(N__37751),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__50006),
            .ce(),
            .sr(N__49111));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2  (
            .in0(N__49470),
            .in1(N__37748),
            .in2(_gnd_net_),
            .in3(N__37733),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__50006),
            .ce(),
            .sr(N__49111));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3  (
            .in0(N__49579),
            .in1(N__39370),
            .in2(_gnd_net_),
            .in3(N__37730),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__50006),
            .ce(),
            .sr(N__49111));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4  (
            .in0(N__49471),
            .in1(N__39396),
            .in2(_gnd_net_),
            .in3(N__37727),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__50006),
            .ce(),
            .sr(N__49111));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5  (
            .in0(N__49580),
            .in1(N__39821),
            .in2(_gnd_net_),
            .in3(N__37961),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__50006),
            .ce(),
            .sr(N__49111));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6  (
            .in0(N__49472),
            .in1(N__39836),
            .in2(_gnd_net_),
            .in3(N__37958),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50006),
            .ce(),
            .sr(N__49111));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_15_9_0  (
            .in0(N__50330),
            .in1(N__42578),
            .in2(_gnd_net_),
            .in3(N__37955),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(N__45115),
            .sr(N__49118));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_15_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_15_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_15_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_15_9_2  (
            .in0(N__50331),
            .in1(N__37935),
            .in2(_gnd_net_),
            .in3(N__42384),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(N__45115),
            .sr(N__49118));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_15_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_15_9_3  (
            .in0(N__37913),
            .in1(N__42520),
            .in2(_gnd_net_),
            .in3(N__50333),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(N__45115),
            .sr(N__49118));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_15_9_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_15_9_4  (
            .in0(N__50328),
            .in1(N__44473),
            .in2(_gnd_net_),
            .in3(N__44512),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(N__45115),
            .sr(N__49118));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_15_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_15_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_15_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_15_9_5  (
            .in0(N__42872),
            .in1(N__50332),
            .in2(_gnd_net_),
            .in3(N__37889),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(N__45115),
            .sr(N__49118));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_15_9_6  (
            .in0(N__50329),
            .in1(N__39575),
            .in2(_gnd_net_),
            .in3(N__43703),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(N__45115),
            .sr(N__49118));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_15_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_15_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_15_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_15_9_7  (
            .in0(N__50520),
            .in1(N__37877),
            .in2(_gnd_net_),
            .in3(N__43983),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49996),
            .ce(N__45115),
            .sr(N__49118));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__38132),
            .in2(N__38171),
            .in3(N__38161),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__38126),
            .in2(N__38108),
            .in3(N__38119),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__38075),
            .in2(N__38099),
            .in3(N__38090),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_10_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_15_10_3  (
            .in0(N__38068),
            .in1(N__38057),
            .in2(N__38051),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__38042),
            .in2(N__38024),
            .in3(N__38035),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_15_10_5  (
            .in0(N__38011),
            .in1(N__38000),
            .in2(N__37994),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_15_10_6  (
            .in0(N__37982),
            .in1(N__37967),
            .in2(N__40193),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__38351),
            .in2(N__38333),
            .in3(N__38344),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__40184),
            .in2(N__38312),
            .in3(N__38323),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__40391),
            .in2(N__38291),
            .in3(N__38302),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__40397),
            .in2(N__38270),
            .in3(N__38281),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__40385),
            .in2(N__38249),
            .in3(N__38260),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__41228),
            .in2(N__38228),
            .in3(N__38239),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_15_11_5  (
            .in0(N__38218),
            .in1(N__38207),
            .in2(N__40094),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__38177),
            .in2(N__38201),
            .in3(N__38188),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__39782),
            .in2(N__39728),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__38429),
            .in2(N__38417),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__40289),
            .in2(N__40343),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__40127),
            .in2(N__40178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__44396),
            .in2(N__44450),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__40082),
            .in2(N__40013),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__39890),
            .in2(N__39956),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__44219),
            .in2(N__44153),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38402),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__44623),
            .in2(N__44648),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__40457),
            .in2(N__40488),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__40379),
            .in2(N__46590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_15_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_15_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__46430),
            .in2(N__38525),
            .in3(N__38501),
            .lcout(\current_shift_inst.un38_control_input_0_s1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_15_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_15_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__40526),
            .in2(N__46591),
            .in3(N__38483),
            .lcout(\current_shift_inst.un38_control_input_0_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_15_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_15_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__46434),
            .in2(N__40373),
            .in3(N__38465),
            .lcout(\current_shift_inst.un38_control_input_0_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__40520),
            .in2(N__46592),
            .in3(N__38450),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__46438),
            .in2(N__40352),
            .in3(N__38432),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__46264),
            .in2(N__38924),
            .in3(N__38612),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__40547),
            .in2(N__46442),
            .in3(N__38597),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__46268),
            .in2(N__41351),
            .in3(N__38582),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__40511),
            .in2(N__46443),
            .in3(N__38567),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__46272),
            .in2(N__41300),
            .in3(N__38552),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__40358),
            .in2(N__46444),
            .in3(N__38537),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__46276),
            .in2(N__41636),
            .in3(N__38534),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__40364),
            .in2(N__46445),
            .in3(N__38531),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__46336),
            .in2(N__39131),
            .in3(N__38528),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__39185),
            .in2(N__46504),
            .in3(N__38741),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__46340),
            .in2(N__39089),
            .in3(N__38738),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__45350),
            .in2(N__46505),
            .in3(N__38720),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__46344),
            .in2(N__39314),
            .in3(N__38702),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__45266),
            .in2(N__46506),
            .in3(N__38687),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__46348),
            .in2(N__38987),
            .in3(N__38672),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__41624),
            .in2(N__46507),
            .in3(N__38654),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__38975),
            .in2(N__46508),
            .in3(N__38639),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__46355),
            .in2(N__39116),
            .in3(N__38831),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__41363),
            .in2(N__46509),
            .in3(N__38828),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__46359),
            .in2(N__39101),
            .in3(N__38825),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__39323),
            .in2(N__46510),
            .in3(N__38807),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__46363),
            .in2(N__38966),
            .in3(N__38789),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_15_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_15_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__40430),
            .in2(N__46511),
            .in3(N__38774),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_15_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_15_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_15_16_7  (
            .in0(N__45999),
            .in1(N__46367),
            .in2(_gnd_net_),
            .in3(N__38771),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_17_0  (
            .in0(N__45986),
            .in1(N__47140),
            .in2(N__46623),
            .in3(N__44598),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_1 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_17_1  (
            .in0(N__46041),
            .in1(N__46524),
            .in2(N__47056),
            .in3(N__45987),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_17_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_17_2  (
            .in0(N__45984),
            .in1(N__46735),
            .in2(N__46622),
            .in3(N__40732),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47049),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_17_4 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_17_4  (
            .in0(N__46525),
            .in1(N__45408),
            .in2(N__46009),
            .in3(N__47012),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_15_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_15_17_5 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_15_17_5  (
            .in0(N__47256),
            .in1(N__45985),
            .in2(N__46700),
            .in3(N__46523),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47255),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46781),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_15_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_15_18_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_15_18_0  (
            .in0(N__41823),
            .in1(N__38912),
            .in2(_gnd_net_),
            .in3(N__38903),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_15_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_15_18_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_15_18_1  (
            .in0(N__38885),
            .in1(N__38876),
            .in2(_gnd_net_),
            .in3(N__41822),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_15_18_2  (
            .in0(N__41826),
            .in1(N__38858),
            .in2(_gnd_net_),
            .in3(N__38849),
            .lcout(\current_shift_inst.control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_18_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_18_3  (
            .in0(N__39074),
            .in1(N__39068),
            .in2(_gnd_net_),
            .in3(N__41824),
            .lcout(\current_shift_inst.control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_15_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_15_18_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_15_18_4  (
            .in0(N__41825),
            .in1(N__39050),
            .in2(_gnd_net_),
            .in3(N__39044),
            .lcout(\current_shift_inst.control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_15_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_15_18_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_15_18_5  (
            .in0(N__41827),
            .in1(N__39023),
            .in2(_gnd_net_),
            .in3(N__39014),
            .lcout(\current_shift_inst.control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_18_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_18_6  (
            .in0(N__45994),
            .in1(N__46527),
            .in2(N__47516),
            .in3(N__45367),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_18_7  (
            .in0(N__46526),
            .in1(N__45995),
            .in2(N__47432),
            .in3(N__45285),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_0  (
            .in0(N__46625),
            .in1(N__45882),
            .in2(N__47384),
            .in3(N__42178),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_19_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_19_1  (
            .in0(N__45883),
            .in1(N__46627),
            .in2(N__48055),
            .in3(N__42052),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_19_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_19_2  (
            .in0(N__46626),
            .in1(N__45887),
            .in2(N__47836),
            .in3(N__41982),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_19_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_19_3  (
            .in0(N__45885),
            .in1(N__46630),
            .in2(N__47969),
            .in3(N__42021),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_4  (
            .in0(N__46628),
            .in1(N__45884),
            .in2(N__48014),
            .in3(N__42080),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_19_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_19_5  (
            .in0(N__45881),
            .in1(N__46629),
            .in2(N__47600),
            .in3(N__45630),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_19_6  (
            .in0(N__46624),
            .in1(N__45886),
            .in2(N__47924),
            .in3(N__41948),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_15_19_7  (
            .in0(N__39167),
            .in1(N__39158),
            .in2(_gnd_net_),
            .in3(N__41862),
            .lcout(\current_shift_inst.control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_20_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_20_0  (
            .in0(N__46637),
            .in1(N__46008),
            .in2(N__47840),
            .in3(N__41983),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_15_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_15_20_1 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_15_20_1  (
            .in0(N__45249),
            .in1(N__46001),
            .in2(N__47648),
            .in3(N__46638),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_2  (
            .in0(N__46002),
            .in1(N__48010),
            .in2(N__46660),
            .in3(N__42079),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_20_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_20_3  (
            .in0(N__46007),
            .in1(N__46632),
            .in2(N__47923),
            .in3(N__41947),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_20_4 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_15_20_4  (
            .in0(N__46631),
            .in1(N__41917),
            .in2(N__47558),
            .in3(N__46005),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_20_5 .LUT_INIT=16'b1111001111110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_20_5  (
            .in0(N__45029),
            .in1(N__46004),
            .in2(N__41012),
            .in3(N__46642),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_20_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_20_6  (
            .in0(N__46003),
            .in1(N__47875),
            .in2(N__46659),
            .in3(N__41716),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_20_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_20_7  (
            .in0(N__46006),
            .in1(N__46636),
            .in2(N__47473),
            .in3(N__45465),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_3_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_3_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_3_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_3_7  (
            .in0(N__40000),
            .in1(N__44059),
            .in2(_gnd_net_),
            .in3(N__50398),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_4_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_4_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_16_4_2  (
            .in0(N__39292),
            .in1(N__42630),
            .in2(_gnd_net_),
            .in3(N__50397),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_4_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_4_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_4_4  (
            .in0(N__39542),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39256),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_4_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_4_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_16_4_6  (
            .in0(N__39541),
            .in1(N__39272),
            .in2(_gnd_net_),
            .in3(N__39255),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_5_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_5_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_16_5_0  (
            .in0(N__39232),
            .in1(N__42666),
            .in2(_gnd_net_),
            .in3(N__50399),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_16_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_16_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_16_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_16_5_1  (
            .in0(_gnd_net_),
            .in1(N__39438),
            .in2(_gnd_net_),
            .in3(N__39469),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_16_5_2  (
            .in0(N__39571),
            .in1(N__43702),
            .in2(_gnd_net_),
            .in3(N__50400),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_16_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_16_5_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_16_5_4  (
            .in0(_gnd_net_),
            .in1(N__39550),
            .in2(_gnd_net_),
            .in3(N__39506),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_5_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39458),
            .in3(N__39437),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_6_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_6_0  (
            .in0(N__39398),
            .in1(N__39376),
            .in2(N__39344),
            .in3(N__39689),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_6_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_6_1  (
            .in0(N__50405),
            .in1(N__40215),
            .in2(_gnd_net_),
            .in3(N__42450),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_16_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_16_6_3 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_16_6_3  (
            .in0(N__39688),
            .in1(N__39397),
            .in2(N__39380),
            .in3(N__39340),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_6_4  (
            .in0(N__43840),
            .in1(N__39874),
            .in2(_gnd_net_),
            .in3(N__50407),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_16_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_16_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_16_6_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_16_6_5  (
            .in0(N__50409),
            .in1(_gnd_net_),
            .in2(N__39347),
            .in3(N__43841),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50037),
            .ce(N__49566),
            .sr(N__49096));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_16_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_16_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_16_6_6  (
            .in0(N__43912),
            .in1(N__39967),
            .in2(_gnd_net_),
            .in3(N__50406),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(elapsed_time_ns_1_RNI69DN9_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_16_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_16_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_16_6_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_16_6_7  (
            .in0(N__50408),
            .in1(_gnd_net_),
            .in2(N__39692),
            .in3(N__43913),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50037),
            .ce(N__49566),
            .sr(N__49096));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_7_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_7_0  (
            .in0(N__39667),
            .in1(N__39648),
            .in2(N__39614),
            .in3(N__39599),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_7_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_16_7_1  (
            .in0(N__39598),
            .in1(N__39666),
            .in2(N__39653),
            .in3(N__39610),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_16_7_2  (
            .in0(N__43251),
            .in1(N__40417),
            .in2(_gnd_net_),
            .in3(N__50291),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(elapsed_time_ns_1_RNI14DN9_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_16_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_16_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_16_7_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_16_7_3  (
            .in0(N__50293),
            .in1(_gnd_net_),
            .in2(N__39617),
            .in3(N__43252),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50030),
            .ce(N__49460),
            .sr(N__49102));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_16_7_4  (
            .in0(N__43308),
            .in1(N__40114),
            .in2(_gnd_net_),
            .in3(N__50290),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(elapsed_time_ns_1_RNI03DN9_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_16_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_16_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_16_7_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_16_7_5  (
            .in0(N__50292),
            .in1(_gnd_net_),
            .in2(N__39602),
            .in3(N__43309),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50030),
            .ce(N__49460),
            .sr(N__49102));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_16_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_16_8_0 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_16_8_0  (
            .in0(N__39845),
            .in1(N__39835),
            .in2(N__50074),
            .in3(N__39820),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_8_1  (
            .in0(N__50556),
            .in1(N__50590),
            .in2(_gnd_net_),
            .in3(N__50281),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_8_3 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_16_8_3  (
            .in0(N__41183),
            .in1(N__41024),
            .in2(N__41141),
            .in3(N__50589),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_8_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__44140),
            .in2(N__39851),
            .in3(N__44101),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(elapsed_time_ns_1_RNIV2EN9_0_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_16_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_16_8_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_16_8_5  (
            .in0(N__44141),
            .in1(_gnd_net_),
            .in2(N__39848),
            .in3(N__50283),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50017),
            .ce(N__49520),
            .sr(N__49107));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_8_6 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_16_8_6  (
            .in0(N__39844),
            .in1(N__39834),
            .in2(N__50075),
            .in3(N__39819),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_16_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_16_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_16_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_16_8_7  (
            .in0(N__41120),
            .in1(N__42977),
            .in2(_gnd_net_),
            .in3(N__50282),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50017),
            .ce(N__49520),
            .sr(N__49107));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_9_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_9_0  (
            .in0(N__39772),
            .in1(N__39751),
            .in2(N__39704),
            .in3(N__39713),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_9_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_9_1  (
            .in0(N__39712),
            .in1(N__39773),
            .in2(N__39752),
            .in3(N__39700),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_16_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_16_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_16_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_16_9_2  (
            .in0(N__40868),
            .in1(N__42812),
            .in2(_gnd_net_),
            .in3(N__50327),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50007),
            .ce(N__45118),
            .sr(N__49112));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_16_9_3  (
            .in0(N__50325),
            .in1(N__42743),
            .in2(_gnd_net_),
            .in3(N__40901),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50007),
            .ce(N__45118),
            .sr(N__49112));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_16_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_16_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_16_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_16_9_4  (
            .in0(N__40843),
            .in1(N__42932),
            .in2(_gnd_net_),
            .in3(N__50326),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50007),
            .ce(N__45118),
            .sr(N__49112));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_16_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_16_10_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_16_10_0  (
            .in0(N__40070),
            .in1(N__40045),
            .in2(N__40037),
            .in3(N__39980),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_16_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_16_10_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_16_10_1  (
            .in0(N__39979),
            .in1(N__40069),
            .in2(N__40049),
            .in3(N__40036),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_16_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_16_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_16_10_2  (
            .in0(N__40001),
            .in1(N__44058),
            .in2(_gnd_net_),
            .in3(N__50511),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49997),
            .ce(N__45116),
            .sr(N__49119));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_16_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_16_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_16_10_4  (
            .in0(N__43911),
            .in1(N__39971),
            .in2(_gnd_net_),
            .in3(N__50512),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49997),
            .ce(N__45116),
            .sr(N__49119));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_16_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_16_10_5 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_16_10_5  (
            .in0(N__39898),
            .in1(N__39944),
            .in2(N__39923),
            .in3(N__39859),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_10_6 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_16_10_6  (
            .in0(N__39943),
            .in1(N__39919),
            .in2(N__39863),
            .in3(N__39899),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_16_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_16_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_16_10_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_16_10_7  (
            .in0(N__50510),
            .in1(N__43839),
            .in2(_gnd_net_),
            .in3(N__39878),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49997),
            .ce(N__45116),
            .sr(N__49119));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_11_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_11_0  (
            .in0(N__40334),
            .in1(N__40309),
            .in2(N__40229),
            .in3(N__40265),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_11_1  (
            .in0(N__40264),
            .in1(N__40333),
            .in2(N__40313),
            .in3(N__40225),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_16_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_16_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_16_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_16_11_2  (
            .in0(N__43427),
            .in1(N__40283),
            .in2(_gnd_net_),
            .in3(N__50354),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(N__45113),
            .sr(N__49126));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_16_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_16_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_16_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_16_11_3  (
            .in0(N__50351),
            .in1(N__40256),
            .in2(_gnd_net_),
            .in3(N__43370),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(N__45113),
            .sr(N__49126));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_16_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_16_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_16_11_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_16_11_6  (
            .in0(N__40217),
            .in1(N__50353),
            .in2(_gnd_net_),
            .in3(N__42454),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(N__45113),
            .sr(N__49126));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_16_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_16_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_16_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_16_11_7  (
            .in0(N__50352),
            .in1(N__41063),
            .in2(_gnd_net_),
            .in3(N__42326),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49986),
            .ce(N__45113),
            .sr(N__49126));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_12_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_16_12_0  (
            .in0(N__40406),
            .in1(N__40103),
            .in2(N__40169),
            .in3(N__40146),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_16_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_16_12_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_16_12_1  (
            .in0(N__40102),
            .in1(N__40168),
            .in2(N__40148),
            .in3(N__40405),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_16_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_16_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_16_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_16_12_2  (
            .in0(N__43313),
            .in1(N__40121),
            .in2(_gnd_net_),
            .in3(N__50509),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49976),
            .ce(N__45111),
            .sr(N__49132));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_16_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_16_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_16_12_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_16_12_3  (
            .in0(N__50507),
            .in1(N__43253),
            .in2(_gnd_net_),
            .in3(N__40421),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49976),
            .ce(N__45111),
            .sr(N__49132));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_16_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_16_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_16_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_16_12_5  (
            .in0(N__50505),
            .in1(N__41174),
            .in2(_gnd_net_),
            .in3(N__43085),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49976),
            .ce(N__45111),
            .sr(N__49132));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_16_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_16_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_16_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_16_12_6  (
            .in0(N__43157),
            .in1(N__41096),
            .in2(_gnd_net_),
            .in3(N__50508),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49976),
            .ce(N__45111),
            .sr(N__49132));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_16_12_7  (
            .in0(N__50506),
            .in1(N__42710),
            .in2(_gnd_net_),
            .in3(N__43028),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49976),
            .ce(N__45111),
            .sr(N__49132));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_13_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_13_0  (
            .in0(N__45911),
            .in1(N__46650),
            .in2(N__46931),
            .in3(N__40609),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_13_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_13_1  (
            .in0(N__46644),
            .in1(N__45913),
            .in2(N__46793),
            .in3(N__44551),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_13_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_13_2  (
            .in0(N__45918),
            .in1(N__46649),
            .in2(N__45215),
            .in3(N__47689),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_13_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_13_3  (
            .in0(N__46648),
            .in1(N__45917),
            .in2(N__47060),
            .in3(N__46045),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_16_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_16_13_4 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_16_13_4  (
            .in0(N__45915),
            .in1(N__46646),
            .in2(N__40709),
            .in3(N__47306),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_13_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_13_5  (
            .in0(N__46643),
            .in1(N__45912),
            .in2(N__46840),
            .in3(N__41338),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_16_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_16_13_6 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_16_13_6  (
            .in0(N__45914),
            .in1(N__46645),
            .in2(N__40736),
            .in3(N__46736),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_13_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_13_7  (
            .in0(N__46647),
            .in1(N__45916),
            .in2(N__47144),
            .in3(N__44605),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_14_0 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_14_0  (
            .in0(N__40489),
            .in1(N__40627),
            .in2(N__40451),
            .in3(N__45826),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48296),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49963),
            .ce(N__47794),
            .sr(N__49145));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40445),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_14_3 .LUT_INIT=16'b1010001110100011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_14_3  (
            .in0(N__40628),
            .in1(N__40450),
            .in2(N__45910),
            .in3(N__40490),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_14_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_14_4  (
            .in0(N__45519),
            .in1(N__40626),
            .in2(_gnd_net_),
            .in3(N__40446),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_16_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_16_14_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_16_14_6  (
            .in0(N__46601),
            .in1(N__45830),
            .in2(N__45028),
            .in3(N__41008),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_16_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_16_15_0 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_16_15_0  (
            .in0(N__47218),
            .in1(N__45991),
            .in2(N__40667),
            .in3(N__46513),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_15_1  (
            .in0(N__45992),
            .in1(N__47219),
            .in2(N__46621),
            .in3(N__40666),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__45993),
            .in2(_gnd_net_),
            .in3(N__46512),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_15_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_15_3  (
            .in0(N__47217),
            .in1(N__45518),
            .in2(_gnd_net_),
            .in3(N__40662),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45671),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_15_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_15_5  (
            .in0(N__45672),
            .in1(_gnd_net_),
            .in2(N__40529),
            .in3(N__45517),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47762),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49954),
            .ce(N__47793),
            .sr(N__49152));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47726),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49954),
            .ce(N__47793),
            .sr(N__49152));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_16_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_16_0  (
            .in0(N__45521),
            .in1(N__46867),
            .in2(_gnd_net_),
            .in3(N__40573),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_16_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_16_1  (
            .in0(N__46827),
            .in1(N__45522),
            .in2(_gnd_net_),
            .in3(N__41331),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_16_2  (
            .in0(N__45525),
            .in1(N__47301),
            .in2(_gnd_net_),
            .in3(N__40695),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_16_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_16_3  (
            .in0(N__46917),
            .in1(N__45520),
            .in2(_gnd_net_),
            .in3(N__40602),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_4  (
            .in0(N__45526),
            .in1(N__47260),
            .in2(_gnd_net_),
            .in3(N__46686),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_16_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_16_5  (
            .in0(N__46731),
            .in1(N__45524),
            .in2(_gnd_net_),
            .in3(N__40728),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_6  (
            .in0(N__45523),
            .in1(N__46782),
            .in2(_gnd_net_),
            .in3(N__44541),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_16_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_16_7  (
            .in0(N__47431),
            .in1(N__45527),
            .in2(_gnd_net_),
            .in3(N__45286),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__40637),
            .in2(N__45085),
            .in3(N__45081),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__41957),
            .in2(_gnd_net_),
            .in3(N__40586),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_17_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42149),
            .in3(N__40562),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__45602),
            .in2(_gnd_net_),
            .in3(N__40748),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__40745),
            .in2(_gnd_net_),
            .in3(N__40739),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__46970),
            .in2(_gnd_net_),
            .in3(N__40712),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__45437),
            .in2(_gnd_net_),
            .in3(N__40679),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__40676),
            .in2(_gnd_net_),
            .in3(N__40670),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__46940),
            .in2(_gnd_net_),
            .in3(N__40649),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__41990),
            .in2(_gnd_net_),
            .in3(N__40646),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__44564),
            .in2(_gnd_net_),
            .in3(N__40643),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__42107),
            .in2(_gnd_net_),
            .in3(N__40640),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__40781),
            .in2(_gnd_net_),
            .in3(N__40775),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(N__46949),
            .in2(_gnd_net_),
            .in3(N__40772),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(N__46958),
            .in2(_gnd_net_),
            .in3(N__40769),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__42260),
            .in2(_gnd_net_),
            .in3(N__40766),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__42137),
            .in2(_gnd_net_),
            .in3(N__40763),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__42245),
            .in2(_gnd_net_),
            .in3(N__40760),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__42227),
            .in2(_gnd_net_),
            .in3(N__40757),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_19_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42131),
            .in3(N__40754),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__42098),
            .in2(_gnd_net_),
            .in3(N__40751),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__42113),
            .in2(_gnd_net_),
            .in3(N__40808),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__42089),
            .in2(_gnd_net_),
            .in3(N__40805),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__42236),
            .in2(_gnd_net_),
            .in3(N__40802),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__42266),
            .in2(_gnd_net_),
            .in3(N__40799),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__42206),
            .in2(_gnd_net_),
            .in3(N__40796),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__42251),
            .in2(_gnd_net_),
            .in3(N__40793),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__42215),
            .in2(_gnd_net_),
            .in3(N__40790),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_20_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42197),
            .in3(N__40787),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40784),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_20_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__46000),
            .in2(_gnd_net_),
            .in3(N__41001),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_17_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_17_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_17_4_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_17_4_6  (
            .in0(N__40860),
            .in1(N__42811),
            .in2(_gnd_net_),
            .in3(N__50501),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50050),
            .ce(N__49550),
            .sr(N__49088));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_5_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_5_0  (
            .in0(N__40973),
            .in1(N__40961),
            .in2(N__40880),
            .in3(N__40936),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_5_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_5_1  (
            .in0(N__40972),
            .in1(N__40960),
            .in2(N__40937),
            .in3(N__40876),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_17_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_17_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_17_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_17_5_2  (
            .in0(N__42741),
            .in1(N__40894),
            .in2(_gnd_net_),
            .in3(N__50403),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(elapsed_time_ns_1_RNI46CN9_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_17_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_17_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_17_5_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_17_5_3  (
            .in0(N__50404),
            .in1(_gnd_net_),
            .in2(N__40883),
            .in3(N__42742),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50047),
            .ce(N__49544),
            .sr(N__49089));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_5_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_5_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_5_4  (
            .in0(N__42804),
            .in1(N__40864),
            .in2(_gnd_net_),
            .in3(N__50402),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_17_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_17_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_17_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_17_5_5  (
            .in0(N__50401),
            .in1(N__40836),
            .in2(_gnd_net_),
            .in3(N__42927),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_17_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_17_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_17_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_17_6_0  (
            .in0(N__40844),
            .in1(N__42928),
            .in2(_gnd_net_),
            .in3(N__50410),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50043),
            .ce(N__49501),
            .sr(N__49093));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_17_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_17_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_17_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_17_6_4  (
            .in0(N__41055),
            .in1(N__42322),
            .in2(_gnd_net_),
            .in3(N__50411),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50043),
            .ce(N__49501),
            .sr(N__49093));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_7_2  (
            .in0(N__43145),
            .in1(N__41089),
            .in2(_gnd_net_),
            .in3(N__50294),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(elapsed_time_ns_1_RNITUBN9_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_3  (
            .in0(N__50296),
            .in1(_gnd_net_),
            .in2(N__41078),
            .in3(N__43146),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50038),
            .ce(N__49563),
            .sr(N__49097));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_7_5  (
            .in0(N__50295),
            .in1(N__41059),
            .in2(_gnd_net_),
            .in3(N__42318),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_17_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_17_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_17_7_7  (
            .in0(N__50297),
            .in1(N__41166),
            .in2(_gnd_net_),
            .in3(N__43078),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50038),
            .ce(N__49563),
            .sr(N__49097));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_17_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_17_8_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(N__42363),
            .in2(_gnd_net_),
            .in3(N__42432),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_17_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_17_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_17_8_2  (
            .in0(N__44505),
            .in1(N__42612),
            .in2(N__43700),
            .in3(N__42648),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_17_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_17_8_3 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__43968),
            .in2(N__41027),
            .in3(N__43905),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_17_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_17_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_17_8_4  (
            .in0(N__43076),
            .in1(N__42317),
            .in2(N__43150),
            .in3(N__43016),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_17_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_17_8_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_17_8_5  (
            .in0(N__42556),
            .in1(N__42503),
            .in2(N__41192),
            .in3(N__41189),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_8_6  (
            .in0(N__43077),
            .in1(N__41170),
            .in2(_gnd_net_),
            .in3(N__50298),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_8_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_8_7  (
            .in0(N__43017),
            .in1(_gnd_net_),
            .in2(N__50420),
            .in3(N__42709),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_17_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_17_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_17_9_0  (
            .in0(N__43476),
            .in1(N__43544),
            .in2(N__43416),
            .in3(N__42726),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_17_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_17_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_17_9_1  (
            .in0(N__42858),
            .in1(N__42917),
            .in2(N__42803),
            .in3(N__42971),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_17_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_17_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_17_9_2  (
            .in0(N__41126),
            .in1(N__41132),
            .in2(N__41150),
            .in3(N__41147),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_17_9_3  (
            .in0(N__44364),
            .in1(N__43236),
            .in2(N__43299),
            .in3(N__43350),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_17_9_4  (
            .in0(N__44139),
            .in1(N__44037),
            .in2(N__44256),
            .in3(N__43827),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_9_5  (
            .in0(N__42972),
            .in1(N__41119),
            .in2(_gnd_net_),
            .in3(N__50302),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(elapsed_time_ns_1_RNI02CN9_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_17_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_17_9_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_17_9_6  (
            .in0(N__50303),
            .in1(_gnd_net_),
            .in2(N__41231),
            .in3(N__42973),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50018),
            .ce(N__45119),
            .sr(N__49108));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0  (
            .in0(N__41535),
            .in1(N__43749),
            .in2(_gnd_net_),
            .in3(N__41216),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__50008),
            .ce(N__41432),
            .sr(N__49113));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1  (
            .in0(N__41541),
            .in1(N__43722),
            .in2(_gnd_net_),
            .in3(N__41213),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__50008),
            .ce(N__41432),
            .sr(N__49113));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2  (
            .in0(N__41536),
            .in1(N__42594),
            .in2(_gnd_net_),
            .in3(N__41210),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__50008),
            .ce(N__41432),
            .sr(N__49113));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3  (
            .in0(N__41542),
            .in1(N__42540),
            .in2(_gnd_net_),
            .in3(N__41207),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__50008),
            .ce(N__41432),
            .sr(N__49113));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4  (
            .in0(N__41537),
            .in1(N__42471),
            .in2(_gnd_net_),
            .in3(N__41204),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__50008),
            .ce(N__41432),
            .sr(N__49113));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5  (
            .in0(N__41543),
            .in1(N__42405),
            .in2(_gnd_net_),
            .in3(N__41201),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__50008),
            .ce(N__41432),
            .sr(N__49113));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6  (
            .in0(N__41538),
            .in1(N__42340),
            .in2(_gnd_net_),
            .in3(N__41198),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__50008),
            .ce(N__41432),
            .sr(N__49113));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7  (
            .in0(N__41544),
            .in1(N__42282),
            .in2(_gnd_net_),
            .in3(N__41195),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__50008),
            .ce(N__41432),
            .sr(N__49113));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0  (
            .in0(N__41560),
            .in1(N__43107),
            .in2(_gnd_net_),
            .in3(N__41258),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__49998),
            .ce(N__41431),
            .sr(N__49120));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1  (
            .in0(N__41548),
            .in1(N__43047),
            .in2(_gnd_net_),
            .in3(N__41255),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__49998),
            .ce(N__41431),
            .sr(N__49120));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2  (
            .in0(N__41557),
            .in1(N__42993),
            .in2(_gnd_net_),
            .in3(N__41252),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__49998),
            .ce(N__41431),
            .sr(N__49120));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3  (
            .in0(N__41545),
            .in1(N__42948),
            .in2(_gnd_net_),
            .in3(N__41249),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__49998),
            .ce(N__41431),
            .sr(N__49120));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4  (
            .in0(N__41558),
            .in1(N__42888),
            .in2(_gnd_net_),
            .in3(N__41246),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__49998),
            .ce(N__41431),
            .sr(N__49120));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5  (
            .in0(N__41546),
            .in1(N__42826),
            .in2(_gnd_net_),
            .in3(N__41243),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__49998),
            .ce(N__41431),
            .sr(N__49120));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6  (
            .in0(N__41559),
            .in1(N__42759),
            .in2(_gnd_net_),
            .in3(N__41240),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__49998),
            .ce(N__41431),
            .sr(N__49120));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7  (
            .in0(N__41547),
            .in1(N__43573),
            .in2(_gnd_net_),
            .in3(N__41237),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__49998),
            .ce(N__41431),
            .sr(N__49120));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0  (
            .in0(N__41549),
            .in1(N__43512),
            .in2(_gnd_net_),
            .in3(N__41234),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__49987),
            .ce(N__41430),
            .sr(N__49127));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1  (
            .in0(N__41561),
            .in1(N__43449),
            .in2(_gnd_net_),
            .in3(N__41285),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__49987),
            .ce(N__41430),
            .sr(N__49127));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2  (
            .in0(N__41550),
            .in1(N__43386),
            .in2(_gnd_net_),
            .in3(N__41282),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__49987),
            .ce(N__41430),
            .sr(N__49127));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3  (
            .in0(N__41562),
            .in1(N__43329),
            .in2(_gnd_net_),
            .in3(N__41279),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__49987),
            .ce(N__41430),
            .sr(N__49127));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4  (
            .in0(N__41551),
            .in1(N__43269),
            .in2(_gnd_net_),
            .in3(N__41276),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__49987),
            .ce(N__41430),
            .sr(N__49127));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5  (
            .in0(N__41563),
            .in1(N__43204),
            .in2(_gnd_net_),
            .in3(N__41273),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__49987),
            .ce(N__41430),
            .sr(N__49127));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6  (
            .in0(N__41552),
            .in1(N__43176),
            .in2(_gnd_net_),
            .in3(N__41270),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__49987),
            .ce(N__41430),
            .sr(N__49127));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7  (
            .in0(N__41564),
            .in1(N__44079),
            .in2(_gnd_net_),
            .in3(N__41267),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__49987),
            .ce(N__41430),
            .sr(N__49127));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0  (
            .in0(N__41553),
            .in1(N__44007),
            .in2(_gnd_net_),
            .in3(N__41264),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__49977),
            .ce(N__41420),
            .sr(N__49133));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1  (
            .in0(N__41539),
            .in1(N__43935),
            .in2(_gnd_net_),
            .in3(N__41261),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__49977),
            .ce(N__41420),
            .sr(N__49133));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2  (
            .in0(N__41554),
            .in1(N__43875),
            .in2(_gnd_net_),
            .in3(N__41573),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__49977),
            .ce(N__41420),
            .sr(N__49133));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3  (
            .in0(N__41540),
            .in1(N__43779),
            .in2(_gnd_net_),
            .in3(N__41570),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__49977),
            .ce(N__41420),
            .sr(N__49133));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4  (
            .in0(N__41555),
            .in1(N__43855),
            .in2(_gnd_net_),
            .in3(N__41567),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__49977),
            .ce(N__41420),
            .sr(N__49133));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5  (
            .in0(N__43804),
            .in1(N__41556),
            .in2(_gnd_net_),
            .in3(N__41435),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49977),
            .ce(N__41420),
            .sr(N__49133));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_0  (
            .in0(N__45838),
            .in1(N__46610),
            .in2(N__45257),
            .in3(N__47644),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_14_1  (
            .in0(N__45909),
            .in1(N__47968),
            .in2(N__46653),
            .in3(N__42026),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_17_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_17_14_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_17_14_2  (
            .in0(N__45835),
            .in1(N__46603),
            .in2(N__47186),
            .in3(N__46094),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_3  (
            .in0(N__46602),
            .in1(N__45834),
            .in2(N__46841),
            .in3(N__41339),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_14_4 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_14_4  (
            .in0(N__47098),
            .in1(N__45907),
            .in2(N__45332),
            .in3(N__46605),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_5  (
            .in0(N__46604),
            .in1(N__45836),
            .in2(N__47102),
            .in3(N__45331),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_17_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_17_14_6 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_17_14_6  (
            .in0(N__45837),
            .in1(N__47011),
            .in2(N__45419),
            .in3(N__46606),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_14_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_17_14_7  (
            .in0(N__45908),
            .in1(N__47341),
            .in2(N__46652),
            .in3(N__45169),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_17_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__45003),
            .in2(N__45055),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_17_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__44973),
            .in2(N__41612),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_17_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__41603),
            .in2(N__44988),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_17_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__44977),
            .in2(N__41597),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_17_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__41588),
            .in2(N__44989),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_17_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__44981),
            .in2(N__41582),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_17_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__41684),
            .in2(N__44990),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_17_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__44985),
            .in2(N__41678),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_17_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__44937),
            .in2(N__41669),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_17_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__44961),
            .in2(N__41660),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_17_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__44934),
            .in2(N__45341),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_17_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__44958),
            .in2(N__44579),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_17_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__44935),
            .in2(N__45302),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_17_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__44959),
            .in2(N__46019),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_17_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__44936),
            .in2(N__45383),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_17_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__44960),
            .in2(N__45428),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_17_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__44918),
            .in2(N__45224),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_17_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__45608),
            .in2(N__44969),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_17_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__44922),
            .in2(N__41900),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_17_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__42122),
            .in2(N__44970),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_17_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__44926),
            .in2(N__45446),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_17_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__41690),
            .in2(N__44971),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_17_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__44930),
            .in2(N__42161),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_17_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__45134),
            .in2(N__44972),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_17_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__44905),
            .in2(N__42035),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_17_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__42062),
            .in2(N__44966),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_17_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__44909),
            .in2(N__41999),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_17_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__41930),
            .in2(N__44967),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_17_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__44913),
            .in2(N__41699),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_17_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__41963),
            .in2(N__44968),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_17_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(N__44917),
            .in2(N__41888),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_18_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_17_18_7  (
            .in0(N__46010),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41876),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_19_0  (
            .in0(N__47868),
            .in1(N__45870),
            .in2(_gnd_net_),
            .in3(N__41715),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_19_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_19_1  (
            .in0(N__45869),
            .in1(N__48003),
            .in2(_gnd_net_),
            .in3(N__42078),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_19_2  (
            .in0(N__48042),
            .in1(N__45588),
            .in2(_gnd_net_),
            .in3(N__42051),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_19_3  (
            .in0(N__47955),
            .in1(N__45872),
            .in2(N__42022),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47163),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_19_5  (
            .in0(N__45871),
            .in1(_gnd_net_),
            .in2(N__41984),
            .in3(N__47823),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46904),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_19_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_19_7  (
            .in0(N__47910),
            .in1(N__45873),
            .in2(_gnd_net_),
            .in3(N__41946),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_20_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_20_0  (
            .in0(N__45585),
            .in1(N__47541),
            .in2(_gnd_net_),
            .in3(N__41916),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_1  (
            .in0(N__47367),
            .in1(N__45586),
            .in2(_gnd_net_),
            .in3(N__42177),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_20_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__46855),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47577),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47446),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_20_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_17_20_5  (
            .in0(N__45587),
            .in1(N__47494),
            .in2(_gnd_net_),
            .in3(N__45366),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47366),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47090),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47408),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47322),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47993),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47624),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47900),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47540),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48033),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47493),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47859),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47945),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47814),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_18_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_18_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_18_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_18_6_2  (
            .in0(N__42705),
            .in1(N__43024),
            .in2(_gnd_net_),
            .in3(N__50521),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50048),
            .ce(N__49564),
            .sr(N__49090));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_7_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_7_0  (
            .in0(_gnd_net_),
            .in1(N__42595),
            .in2(N__43757),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_18_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50044),
            .ce(N__43652),
            .sr(N__49094));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_7_1  (
            .in0(_gnd_net_),
            .in1(N__42541),
            .in2(N__43730),
            .in3(N__42599),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50044),
            .ce(N__43652),
            .sr(N__49094));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_7_2  (
            .in0(_gnd_net_),
            .in1(N__42596),
            .in2(N__42478),
            .in3(N__42545),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50044),
            .ce(N__43652),
            .sr(N__49094));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_7_3  (
            .in0(_gnd_net_),
            .in1(N__42542),
            .in2(N__42412),
            .in3(N__42482),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50044),
            .ce(N__43652),
            .sr(N__49094));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_7_4  (
            .in0(_gnd_net_),
            .in1(N__42346),
            .in2(N__42479),
            .in3(N__42416),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50044),
            .ce(N__43652),
            .sr(N__49094));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_7_5  (
            .in0(_gnd_net_),
            .in1(N__42289),
            .in2(N__42413),
            .in3(N__42350),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50044),
            .ce(N__43652),
            .sr(N__49094));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_7_6  (
            .in0(_gnd_net_),
            .in1(N__42347),
            .in2(N__43120),
            .in3(N__42296),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50044),
            .ce(N__43652),
            .sr(N__49094));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_7_7  (
            .in0(_gnd_net_),
            .in1(N__43054),
            .in2(N__42293),
            .in3(N__43124),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50044),
            .ce(N__43652),
            .sr(N__49094));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_8_0  (
            .in0(_gnd_net_),
            .in1(N__42994),
            .in2(N__43121),
            .in3(N__43058),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_18_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50039),
            .ce(N__43651),
            .sr(N__49098));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(N__42949),
            .in2(N__43055),
            .in3(N__42998),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50039),
            .ce(N__43651),
            .sr(N__49098));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_8_2  (
            .in0(_gnd_net_),
            .in1(N__42995),
            .in2(N__42895),
            .in3(N__42953),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50039),
            .ce(N__43651),
            .sr(N__49098));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(N__42950),
            .in2(N__42838),
            .in3(N__42899),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50039),
            .ce(N__43651),
            .sr(N__49098));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(N__42766),
            .in2(N__42896),
            .in3(N__42842),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50039),
            .ce(N__43651),
            .sr(N__49098));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(N__43579),
            .in2(N__42839),
            .in3(N__42773),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50039),
            .ce(N__43651),
            .sr(N__49098));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_8_6  (
            .in0(_gnd_net_),
            .in1(N__43519),
            .in2(N__42770),
            .in3(N__42713),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50039),
            .ce(N__43651),
            .sr(N__49098));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_8_7  (
            .in0(_gnd_net_),
            .in1(N__43580),
            .in2(N__43460),
            .in3(N__43526),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50039),
            .ce(N__43651),
            .sr(N__49098));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_9_0  (
            .in0(_gnd_net_),
            .in1(N__43387),
            .in2(N__43523),
            .in3(N__43463),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50031),
            .ce(N__43650),
            .sr(N__49103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_9_1  (
            .in0(_gnd_net_),
            .in1(N__43330),
            .in2(N__43459),
            .in3(N__43391),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50031),
            .ce(N__43650),
            .sr(N__49103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(N__43388),
            .in2(N__43276),
            .in3(N__43334),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50031),
            .ce(N__43650),
            .sr(N__49103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_9_3  (
            .in0(_gnd_net_),
            .in1(N__43331),
            .in2(N__43216),
            .in3(N__43280),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50031),
            .ce(N__43650),
            .sr(N__49103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_9_4  (
            .in0(_gnd_net_),
            .in1(N__43183),
            .in2(N__43277),
            .in3(N__43220),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50031),
            .ce(N__43650),
            .sr(N__49103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_9_5  (
            .in0(_gnd_net_),
            .in1(N__44086),
            .in2(N__43217),
            .in3(N__43190),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50031),
            .ce(N__43650),
            .sr(N__49103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_9_6  (
            .in0(_gnd_net_),
            .in1(N__44014),
            .in2(N__43187),
            .in3(N__43160),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50031),
            .ce(N__43650),
            .sr(N__49103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_9_7  (
            .in0(_gnd_net_),
            .in1(N__43942),
            .in2(N__44090),
            .in3(N__44021),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50031),
            .ce(N__43650),
            .sr(N__49103));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__43876),
            .in2(N__44018),
            .in3(N__43946),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50019),
            .ce(N__43649),
            .sr(N__49109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(N__43786),
            .in2(N__43943),
            .in3(N__43880),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50019),
            .ce(N__43649),
            .sr(N__49109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(N__43877),
            .in2(N__43859),
            .in3(N__43811),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50019),
            .ce(N__43649),
            .sr(N__49109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(N__43808),
            .in2(N__43790),
            .in3(N__43763),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50019),
            .ce(N__43649),
            .sr(N__49109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43760),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50019),
            .ce(N__43649),
            .sr(N__49109));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43750),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50009),
            .ce(N__43645),
            .sr(N__49114));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43723),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50009),
            .ce(N__43645),
            .sr(N__49114));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_4  (
            .in0(N__44466),
            .in1(N__44499),
            .in2(_gnd_net_),
            .in3(N__50469),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_12_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_12_0  (
            .in0(N__44437),
            .in1(N__44416),
            .in2(N__44231),
            .in3(N__44321),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_12_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_12_1  (
            .in0(N__44320),
            .in1(N__44438),
            .in2(N__44420),
            .in3(N__44227),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_18_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_18_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_18_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_18_12_2  (
            .in0(N__44385),
            .in1(N__44351),
            .in2(_gnd_net_),
            .in3(N__50514),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49999),
            .ce(N__45117),
            .sr(N__49121));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_18_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_18_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_18_12_3  (
            .in0(N__50513),
            .in1(N__44312),
            .in2(_gnd_net_),
            .in3(N__44271),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49999),
            .ce(N__45117),
            .sr(N__49121));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_18_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_18_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_18_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_18_12_4  (
            .in0(N__50588),
            .in1(N__50558),
            .in2(_gnd_net_),
            .in3(N__50515),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49999),
            .ce(N__45117),
            .sr(N__49121));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_12_5 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_12_5  (
            .in0(N__45127),
            .in1(N__44200),
            .in2(N__44177),
            .in3(N__44209),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_18_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_18_12_6 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_18_12_6  (
            .in0(N__44210),
            .in1(N__45128),
            .in2(N__44201),
            .in3(N__44176),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_18_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_18_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_18_13_6  (
            .in0(N__44138),
            .in1(N__44111),
            .in2(_gnd_net_),
            .in3(N__50528),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49988),
            .ce(N__45114),
            .sr(N__49128));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45086),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_14_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__45813),
            .in2(N__45059),
            .in3(N__45685),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47757),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49978),
            .ce(N__47795),
            .sr(N__49134));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_18_14_4  (
            .in0(N__45056),
            .in1(N__44986),
            .in2(_gnd_net_),
            .in3(N__45035),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_18_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_18_14_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_18_14_5  (
            .in0(N__44987),
            .in1(_gnd_net_),
            .in2(N__44651),
            .in3(N__44641),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_14_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_18_14_6  (
            .in0(N__47130),
            .in1(N__45572),
            .in2(_gnd_net_),
            .in3(N__44606),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47129),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_18_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_18_15_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_18_15_0  (
            .in0(N__46587),
            .in1(N__45960),
            .in2(N__46789),
            .in3(N__44552),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_15_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_18_15_1  (
            .in0(N__47685),
            .in1(N__45552),
            .in2(_gnd_net_),
            .in3(N__45210),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_18_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_18_15_2 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_18_15_2  (
            .in0(N__45551),
            .in1(N__47007),
            .in2(N__45415),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_4  (
            .in0(N__46589),
            .in1(N__45961),
            .in2(N__47512),
            .in3(N__45374),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_15_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_18_15_5  (
            .in0(N__47179),
            .in1(N__45549),
            .in2(_gnd_net_),
            .in3(N__46092),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_15_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_18_15_6  (
            .in0(N__45550),
            .in1(N__47091),
            .in2(_gnd_net_),
            .in3(N__45327),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_15_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_18_15_7  (
            .in0(N__45962),
            .in1(N__46588),
            .in2(N__45293),
            .in3(N__47421),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_16_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_18_16_0  (
            .in0(N__47643),
            .in1(N__45590),
            .in2(_gnd_net_),
            .in3(N__45250),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_18_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_18_16_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_18_16_1  (
            .in0(N__45959),
            .in1(N__46658),
            .in2(N__47690),
            .in3(N__45211),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_18_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_18_16_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_18_16_2  (
            .in0(N__47340),
            .in1(N__45591),
            .in2(_gnd_net_),
            .in3(N__45168),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_18_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_18_16_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_18_16_3  (
            .in0(N__45957),
            .in1(N__46657),
            .in2(N__47261),
            .in3(N__46699),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_18_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_18_16_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_18_16_4  (
            .in0(N__47178),
            .in1(N__45958),
            .in2(N__46661),
            .in3(N__46093),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_16_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_18_16_6  (
            .in0(N__47048),
            .in1(N__45589),
            .in2(_gnd_net_),
            .in3(N__46046),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_18_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_18_16_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_18_16_7  (
            .in0(N__45956),
            .in1(N__45695),
            .in2(_gnd_net_),
            .in3(N__45686),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_18_17_0  (
            .in0(N__45592),
            .in1(N__47595),
            .in2(_gnd_net_),
            .in3(N__45637),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46818),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_18_17_4  (
            .in0(N__45593),
            .in1(N__47460),
            .in2(_gnd_net_),
            .in3(N__45472),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47283),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46714),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47675),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47003),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47200),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__48253),
            .in2(N__47722),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49940),
            .ce(N__47791),
            .sr(N__49162));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__48232),
            .in2(N__48292),
            .in3(N__46844),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49940),
            .ce(N__47791),
            .sr(N__49162));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__48254),
            .in2(N__48212),
            .in3(N__46796),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49940),
            .ce(N__47791),
            .sr(N__49162));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__48233),
            .in2(N__48182),
            .in3(N__46739),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49940),
            .ce(N__47791),
            .sr(N__49162));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__48211),
            .in2(N__48151),
            .in3(N__46703),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49940),
            .ce(N__47791),
            .sr(N__49162));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__48181),
            .in2(N__48121),
            .in3(N__47264),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49940),
            .ce(N__47791),
            .sr(N__49162));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__48088),
            .in2(N__48152),
            .in3(N__47222),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49940),
            .ce(N__47791),
            .sr(N__49162));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__48544),
            .in2(N__48122),
            .in3(N__47189),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49940),
            .ce(N__47791),
            .sr(N__49162));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__48517),
            .in2(N__48092),
            .in3(N__47147),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49933),
            .ce(N__47790),
            .sr(N__49167));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__48493),
            .in2(N__48548),
            .in3(N__47105),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49933),
            .ce(N__47790),
            .sr(N__49167));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__48518),
            .in2(N__48469),
            .in3(N__47063),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49933),
            .ce(N__47790),
            .sr(N__49167));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__48494),
            .in2(N__48439),
            .in3(N__47015),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49933),
            .ce(N__47790),
            .sr(N__49167));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__48409),
            .in2(N__48470),
            .in3(N__46973),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49933),
            .ce(N__47790),
            .sr(N__49167));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__48382),
            .in2(N__48440),
            .in3(N__47651),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49933),
            .ce(N__47790),
            .sr(N__49167));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__48410),
            .in2(N__48355),
            .in3(N__47603),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49933),
            .ce(N__47790),
            .sr(N__49167));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(N__48322),
            .in2(N__48386),
            .in3(N__47561),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49933),
            .ce(N__47790),
            .sr(N__49167));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__48760),
            .in2(N__48356),
            .in3(N__47519),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49927),
            .ce(N__47789),
            .sr(N__49172));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__48323),
            .in2(N__48739),
            .in3(N__47477),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49927),
            .ce(N__47789),
            .sr(N__49172));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__48761),
            .in2(N__48713),
            .in3(N__47435),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49927),
            .ce(N__47789),
            .sr(N__49172));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(N__48682),
            .in2(N__48740),
            .in3(N__47387),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49927),
            .ce(N__47789),
            .sr(N__49172));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_21_4  (
            .in0(_gnd_net_),
            .in1(N__48712),
            .in2(N__48658),
            .in3(N__47348),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49927),
            .ce(N__47789),
            .sr(N__49172));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_21_5  (
            .in0(_gnd_net_),
            .in1(N__48628),
            .in2(N__48686),
            .in3(N__48062),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49927),
            .ce(N__47789),
            .sr(N__49172));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_21_6  (
            .in0(_gnd_net_),
            .in1(N__48604),
            .in2(N__48659),
            .in3(N__48017),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49927),
            .ce(N__47789),
            .sr(N__49172));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(N__48629),
            .in2(N__48578),
            .in3(N__47972),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49927),
            .ce(N__47789),
            .sr(N__49172));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(N__50851),
            .in2(N__48608),
            .in3(N__47927),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_18_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49922),
            .ce(N__47788),
            .sr(N__49178));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__48577),
            .in2(N__50827),
            .in3(N__47879),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49922),
            .ce(N__47788),
            .sr(N__49178));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__50801),
            .in2(N__50855),
            .in3(N__47843),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49922),
            .ce(N__47788),
            .sr(N__49178));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(N__50657),
            .in2(N__50828),
            .in3(N__47798),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49922),
            .ce(N__47788),
            .sr(N__49178));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47765),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_18_23_0  (
            .in0(N__50758),
            .in1(N__47712),
            .in2(_gnd_net_),
            .in3(N__47693),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_23_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__49915),
            .ce(N__50633),
            .sr(N__49182));
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_18_23_1  (
            .in0(N__50754),
            .in1(N__48276),
            .in2(_gnd_net_),
            .in3(N__48257),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__49915),
            .ce(N__50633),
            .sr(N__49182));
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_18_23_2  (
            .in0(N__50759),
            .in1(N__48252),
            .in2(_gnd_net_),
            .in3(N__48236),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__49915),
            .ce(N__50633),
            .sr(N__49182));
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_18_23_3  (
            .in0(N__50755),
            .in1(N__48231),
            .in2(_gnd_net_),
            .in3(N__48215),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__49915),
            .ce(N__50633),
            .sr(N__49182));
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_18_23_4  (
            .in0(N__50760),
            .in1(N__48201),
            .in2(_gnd_net_),
            .in3(N__48185),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__49915),
            .ce(N__50633),
            .sr(N__49182));
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_18_23_5  (
            .in0(N__50756),
            .in1(N__48171),
            .in2(_gnd_net_),
            .in3(N__48155),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__49915),
            .ce(N__50633),
            .sr(N__49182));
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_18_23_6  (
            .in0(N__50761),
            .in1(N__48139),
            .in2(_gnd_net_),
            .in3(N__48125),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__49915),
            .ce(N__50633),
            .sr(N__49182));
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_18_23_7  (
            .in0(N__50757),
            .in1(N__48109),
            .in2(_gnd_net_),
            .in3(N__48095),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__49915),
            .ce(N__50633),
            .sr(N__49182));
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_18_24_0  (
            .in0(N__50779),
            .in1(N__48081),
            .in2(_gnd_net_),
            .in3(N__48065),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__49911),
            .ce(N__50641),
            .sr(N__49188));
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_18_24_1  (
            .in0(N__50783),
            .in1(N__48537),
            .in2(_gnd_net_),
            .in3(N__48521),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__49911),
            .ce(N__50641),
            .sr(N__49188));
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_18_24_2  (
            .in0(N__50776),
            .in1(N__48511),
            .in2(_gnd_net_),
            .in3(N__48497),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__49911),
            .ce(N__50641),
            .sr(N__49188));
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_18_24_3  (
            .in0(N__50780),
            .in1(N__48487),
            .in2(_gnd_net_),
            .in3(N__48473),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__49911),
            .ce(N__50641),
            .sr(N__49188));
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_18_24_4  (
            .in0(N__50777),
            .in1(N__48457),
            .in2(_gnd_net_),
            .in3(N__48443),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__49911),
            .ce(N__50641),
            .sr(N__49188));
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_18_24_5  (
            .in0(N__50781),
            .in1(N__48427),
            .in2(_gnd_net_),
            .in3(N__48413),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__49911),
            .ce(N__50641),
            .sr(N__49188));
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_18_24_6  (
            .in0(N__50778),
            .in1(N__48403),
            .in2(_gnd_net_),
            .in3(N__48389),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__49911),
            .ce(N__50641),
            .sr(N__49188));
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_18_24_7  (
            .in0(N__50782),
            .in1(N__48375),
            .in2(_gnd_net_),
            .in3(N__48359),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__49911),
            .ce(N__50641),
            .sr(N__49188));
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_18_25_0  (
            .in0(N__50762),
            .in1(N__48342),
            .in2(_gnd_net_),
            .in3(N__48326),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_25_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__49908),
            .ce(N__50640),
            .sr(N__49193));
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_18_25_1  (
            .in0(N__50770),
            .in1(N__48315),
            .in2(_gnd_net_),
            .in3(N__48299),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__49908),
            .ce(N__50640),
            .sr(N__49193));
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_18_25_2  (
            .in0(N__50763),
            .in1(N__48759),
            .in2(_gnd_net_),
            .in3(N__48743),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__49908),
            .ce(N__50640),
            .sr(N__49193));
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_18_25_3  (
            .in0(N__50771),
            .in1(N__48732),
            .in2(_gnd_net_),
            .in3(N__48716),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__49908),
            .ce(N__50640),
            .sr(N__49193));
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_18_25_4  (
            .in0(N__50764),
            .in1(N__48708),
            .in2(_gnd_net_),
            .in3(N__48689),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__49908),
            .ce(N__50640),
            .sr(N__49193));
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_25_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_18_25_5  (
            .in0(N__50772),
            .in1(N__48681),
            .in2(_gnd_net_),
            .in3(N__48662),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__49908),
            .ce(N__50640),
            .sr(N__49193));
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_25_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_18_25_6  (
            .in0(N__50765),
            .in1(N__48646),
            .in2(_gnd_net_),
            .in3(N__48632),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__49908),
            .ce(N__50640),
            .sr(N__49193));
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_25_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_18_25_7  (
            .in0(N__50773),
            .in1(N__48627),
            .in2(_gnd_net_),
            .in3(N__48611),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__49908),
            .ce(N__50640),
            .sr(N__49193));
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_26_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_18_26_0  (
            .in0(N__50766),
            .in1(N__48597),
            .in2(_gnd_net_),
            .in3(N__48581),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_18_26_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__49905),
            .ce(N__50642),
            .sr(N__49199));
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_26_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_26_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_18_26_1  (
            .in0(N__50774),
            .in1(N__48567),
            .in2(_gnd_net_),
            .in3(N__48551),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__49905),
            .ce(N__50642),
            .sr(N__49199));
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_26_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_18_26_2  (
            .in0(N__50767),
            .in1(N__50850),
            .in2(_gnd_net_),
            .in3(N__50831),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__49905),
            .ce(N__50642),
            .sr(N__49199));
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_26_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_18_26_3  (
            .in0(N__50775),
            .in1(N__50820),
            .in2(_gnd_net_),
            .in3(N__50804),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__49905),
            .ce(N__50642),
            .sr(N__49199));
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_26_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_26_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_18_26_4  (
            .in0(N__50768),
            .in1(N__50800),
            .in2(_gnd_net_),
            .in3(N__50786),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__49905),
            .ce(N__50642),
            .sr(N__49199));
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_26_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_26_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_18_26_5  (
            .in0(N__50656),
            .in1(N__50769),
            .in2(_gnd_net_),
            .in3(N__50660),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49905),
            .ce(N__50642),
            .sr(N__49199));
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_2.C_ON=1'b0;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_2 (
            .in0(N__50054),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clock_output_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_20_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_20_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_20_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_20_9_4  (
            .in0(N__50591),
            .in1(N__50557),
            .in2(_gnd_net_),
            .in3(N__50524),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50045),
            .ce(N__49542),
            .sr(N__49104));
endmodule // MAIN
