// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Nov 15 2024 21:13:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    error_pin,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    input error_pin;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__50511;
    wire N__50510;
    wire N__50509;
    wire N__50500;
    wire N__50499;
    wire N__50498;
    wire N__50491;
    wire N__50490;
    wire N__50489;
    wire N__50482;
    wire N__50481;
    wire N__50480;
    wire N__50473;
    wire N__50472;
    wire N__50471;
    wire N__50464;
    wire N__50463;
    wire N__50462;
    wire N__50455;
    wire N__50454;
    wire N__50453;
    wire N__50446;
    wire N__50445;
    wire N__50444;
    wire N__50437;
    wire N__50436;
    wire N__50435;
    wire N__50428;
    wire N__50427;
    wire N__50426;
    wire N__50419;
    wire N__50418;
    wire N__50417;
    wire N__50410;
    wire N__50409;
    wire N__50408;
    wire N__50401;
    wire N__50400;
    wire N__50399;
    wire N__50382;
    wire N__50379;
    wire N__50376;
    wire N__50375;
    wire N__50372;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50362;
    wire N__50355;
    wire N__50352;
    wire N__50351;
    wire N__50348;
    wire N__50345;
    wire N__50344;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50325;
    wire N__50324;
    wire N__50323;
    wire N__50320;
    wire N__50319;
    wire N__50316;
    wire N__50313;
    wire N__50310;
    wire N__50307;
    wire N__50304;
    wire N__50301;
    wire N__50296;
    wire N__50293;
    wire N__50288;
    wire N__50283;
    wire N__50280;
    wire N__50279;
    wire N__50278;
    wire N__50277;
    wire N__50274;
    wire N__50271;
    wire N__50268;
    wire N__50265;
    wire N__50260;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50238;
    wire N__50235;
    wire N__50234;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50226;
    wire N__50223;
    wire N__50218;
    wire N__50215;
    wire N__50214;
    wire N__50211;
    wire N__50208;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50196;
    wire N__50191;
    wire N__50184;
    wire N__50183;
    wire N__50182;
    wire N__50181;
    wire N__50180;
    wire N__50179;
    wire N__50178;
    wire N__50177;
    wire N__50176;
    wire N__50175;
    wire N__50174;
    wire N__50173;
    wire N__50172;
    wire N__50171;
    wire N__50170;
    wire N__50169;
    wire N__50168;
    wire N__50167;
    wire N__50166;
    wire N__50165;
    wire N__50164;
    wire N__50163;
    wire N__50162;
    wire N__50161;
    wire N__50160;
    wire N__50159;
    wire N__50150;
    wire N__50149;
    wire N__50148;
    wire N__50147;
    wire N__50146;
    wire N__50137;
    wire N__50128;
    wire N__50123;
    wire N__50114;
    wire N__50105;
    wire N__50096;
    wire N__50093;
    wire N__50084;
    wire N__50079;
    wire N__50076;
    wire N__50073;
    wire N__50068;
    wire N__50063;
    wire N__50060;
    wire N__50055;
    wire N__50052;
    wire N__50043;
    wire N__50042;
    wire N__50039;
    wire N__50036;
    wire N__50035;
    wire N__50032;
    wire N__50027;
    wire N__50022;
    wire N__50019;
    wire N__50016;
    wire N__50013;
    wire N__50010;
    wire N__50007;
    wire N__50006;
    wire N__50003;
    wire N__50000;
    wire N__49995;
    wire N__49992;
    wire N__49991;
    wire N__49990;
    wire N__49987;
    wire N__49982;
    wire N__49979;
    wire N__49974;
    wire N__49973;
    wire N__49972;
    wire N__49971;
    wire N__49968;
    wire N__49961;
    wire N__49956;
    wire N__49955;
    wire N__49954;
    wire N__49953;
    wire N__49952;
    wire N__49951;
    wire N__49950;
    wire N__49949;
    wire N__49948;
    wire N__49947;
    wire N__49946;
    wire N__49945;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49941;
    wire N__49940;
    wire N__49939;
    wire N__49938;
    wire N__49937;
    wire N__49936;
    wire N__49935;
    wire N__49934;
    wire N__49933;
    wire N__49932;
    wire N__49931;
    wire N__49930;
    wire N__49929;
    wire N__49928;
    wire N__49927;
    wire N__49926;
    wire N__49925;
    wire N__49924;
    wire N__49923;
    wire N__49922;
    wire N__49921;
    wire N__49920;
    wire N__49919;
    wire N__49918;
    wire N__49917;
    wire N__49916;
    wire N__49915;
    wire N__49914;
    wire N__49913;
    wire N__49912;
    wire N__49911;
    wire N__49910;
    wire N__49909;
    wire N__49908;
    wire N__49907;
    wire N__49906;
    wire N__49905;
    wire N__49904;
    wire N__49903;
    wire N__49902;
    wire N__49901;
    wire N__49900;
    wire N__49899;
    wire N__49898;
    wire N__49897;
    wire N__49896;
    wire N__49895;
    wire N__49894;
    wire N__49893;
    wire N__49892;
    wire N__49891;
    wire N__49890;
    wire N__49889;
    wire N__49888;
    wire N__49887;
    wire N__49886;
    wire N__49885;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49881;
    wire N__49880;
    wire N__49879;
    wire N__49878;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49874;
    wire N__49873;
    wire N__49872;
    wire N__49871;
    wire N__49870;
    wire N__49869;
    wire N__49868;
    wire N__49867;
    wire N__49866;
    wire N__49865;
    wire N__49864;
    wire N__49863;
    wire N__49862;
    wire N__49861;
    wire N__49860;
    wire N__49859;
    wire N__49858;
    wire N__49857;
    wire N__49856;
    wire N__49855;
    wire N__49854;
    wire N__49853;
    wire N__49852;
    wire N__49851;
    wire N__49850;
    wire N__49849;
    wire N__49848;
    wire N__49847;
    wire N__49846;
    wire N__49845;
    wire N__49844;
    wire N__49843;
    wire N__49842;
    wire N__49841;
    wire N__49840;
    wire N__49839;
    wire N__49838;
    wire N__49837;
    wire N__49836;
    wire N__49835;
    wire N__49834;
    wire N__49833;
    wire N__49832;
    wire N__49831;
    wire N__49830;
    wire N__49829;
    wire N__49828;
    wire N__49827;
    wire N__49826;
    wire N__49825;
    wire N__49824;
    wire N__49823;
    wire N__49822;
    wire N__49821;
    wire N__49820;
    wire N__49819;
    wire N__49818;
    wire N__49817;
    wire N__49816;
    wire N__49815;
    wire N__49814;
    wire N__49813;
    wire N__49812;
    wire N__49811;
    wire N__49810;
    wire N__49809;
    wire N__49808;
    wire N__49807;
    wire N__49806;
    wire N__49805;
    wire N__49804;
    wire N__49803;
    wire N__49802;
    wire N__49801;
    wire N__49800;
    wire N__49799;
    wire N__49482;
    wire N__49479;
    wire N__49478;
    wire N__49477;
    wire N__49476;
    wire N__49473;
    wire N__49470;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49458;
    wire N__49455;
    wire N__49454;
    wire N__49453;
    wire N__49452;
    wire N__49451;
    wire N__49450;
    wire N__49447;
    wire N__49446;
    wire N__49445;
    wire N__49444;
    wire N__49443;
    wire N__49442;
    wire N__49441;
    wire N__49440;
    wire N__49439;
    wire N__49438;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49431;
    wire N__49430;
    wire N__49429;
    wire N__49428;
    wire N__49427;
    wire N__49426;
    wire N__49425;
    wire N__49424;
    wire N__49423;
    wire N__49422;
    wire N__49421;
    wire N__49420;
    wire N__49419;
    wire N__49418;
    wire N__49417;
    wire N__49416;
    wire N__49415;
    wire N__49414;
    wire N__49413;
    wire N__49412;
    wire N__49411;
    wire N__49410;
    wire N__49409;
    wire N__49408;
    wire N__49407;
    wire N__49406;
    wire N__49405;
    wire N__49404;
    wire N__49403;
    wire N__49402;
    wire N__49401;
    wire N__49400;
    wire N__49399;
    wire N__49398;
    wire N__49397;
    wire N__49396;
    wire N__49395;
    wire N__49394;
    wire N__49393;
    wire N__49392;
    wire N__49391;
    wire N__49390;
    wire N__49389;
    wire N__49388;
    wire N__49387;
    wire N__49386;
    wire N__49385;
    wire N__49384;
    wire N__49383;
    wire N__49382;
    wire N__49381;
    wire N__49380;
    wire N__49379;
    wire N__49378;
    wire N__49377;
    wire N__49376;
    wire N__49375;
    wire N__49374;
    wire N__49373;
    wire N__49372;
    wire N__49371;
    wire N__49370;
    wire N__49369;
    wire N__49368;
    wire N__49367;
    wire N__49366;
    wire N__49365;
    wire N__49364;
    wire N__49363;
    wire N__49362;
    wire N__49361;
    wire N__49360;
    wire N__49359;
    wire N__49358;
    wire N__49357;
    wire N__49356;
    wire N__49355;
    wire N__49354;
    wire N__49353;
    wire N__49352;
    wire N__49351;
    wire N__49350;
    wire N__49349;
    wire N__49348;
    wire N__49347;
    wire N__49346;
    wire N__49345;
    wire N__49344;
    wire N__49343;
    wire N__49342;
    wire N__49341;
    wire N__49340;
    wire N__49339;
    wire N__49338;
    wire N__49337;
    wire N__49336;
    wire N__49335;
    wire N__49334;
    wire N__49333;
    wire N__49332;
    wire N__49331;
    wire N__49330;
    wire N__49329;
    wire N__49328;
    wire N__49327;
    wire N__49326;
    wire N__49325;
    wire N__49324;
    wire N__49323;
    wire N__49322;
    wire N__49321;
    wire N__49320;
    wire N__49319;
    wire N__49318;
    wire N__49317;
    wire N__49316;
    wire N__49315;
    wire N__49314;
    wire N__49313;
    wire N__49312;
    wire N__49311;
    wire N__49310;
    wire N__49309;
    wire N__49308;
    wire N__49307;
    wire N__49306;
    wire N__49305;
    wire N__49304;
    wire N__49303;
    wire N__49302;
    wire N__49301;
    wire N__49300;
    wire N__49299;
    wire N__49298;
    wire N__49297;
    wire N__49296;
    wire N__49295;
    wire N__49294;
    wire N__49293;
    wire N__49292;
    wire N__49291;
    wire N__48960;
    wire N__48957;
    wire N__48954;
    wire N__48953;
    wire N__48952;
    wire N__48951;
    wire N__48948;
    wire N__48945;
    wire N__48944;
    wire N__48941;
    wire N__48940;
    wire N__48937;
    wire N__48936;
    wire N__48933;
    wire N__48932;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48910;
    wire N__48905;
    wire N__48902;
    wire N__48899;
    wire N__48896;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48882;
    wire N__48881;
    wire N__48878;
    wire N__48875;
    wire N__48870;
    wire N__48869;
    wire N__48868;
    wire N__48867;
    wire N__48866;
    wire N__48865;
    wire N__48864;
    wire N__48863;
    wire N__48862;
    wire N__48861;
    wire N__48860;
    wire N__48859;
    wire N__48858;
    wire N__48857;
    wire N__48856;
    wire N__48855;
    wire N__48854;
    wire N__48853;
    wire N__48852;
    wire N__48851;
    wire N__48850;
    wire N__48849;
    wire N__48846;
    wire N__48843;
    wire N__48840;
    wire N__48839;
    wire N__48838;
    wire N__48837;
    wire N__48836;
    wire N__48835;
    wire N__48818;
    wire N__48803;
    wire N__48800;
    wire N__48797;
    wire N__48796;
    wire N__48793;
    wire N__48790;
    wire N__48785;
    wire N__48782;
    wire N__48781;
    wire N__48780;
    wire N__48775;
    wire N__48768;
    wire N__48763;
    wire N__48758;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48734;
    wire N__48731;
    wire N__48730;
    wire N__48729;
    wire N__48722;
    wire N__48719;
    wire N__48716;
    wire N__48713;
    wire N__48710;
    wire N__48707;
    wire N__48704;
    wire N__48701;
    wire N__48696;
    wire N__48689;
    wire N__48686;
    wire N__48683;
    wire N__48680;
    wire N__48677;
    wire N__48672;
    wire N__48663;
    wire N__48660;
    wire N__48657;
    wire N__48654;
    wire N__48651;
    wire N__48648;
    wire N__48647;
    wire N__48646;
    wire N__48645;
    wire N__48644;
    wire N__48643;
    wire N__48642;
    wire N__48641;
    wire N__48640;
    wire N__48639;
    wire N__48638;
    wire N__48629;
    wire N__48628;
    wire N__48627;
    wire N__48626;
    wire N__48625;
    wire N__48624;
    wire N__48623;
    wire N__48622;
    wire N__48619;
    wire N__48612;
    wire N__48607;
    wire N__48604;
    wire N__48601;
    wire N__48592;
    wire N__48585;
    wire N__48584;
    wire N__48583;
    wire N__48582;
    wire N__48581;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48563;
    wire N__48552;
    wire N__48551;
    wire N__48550;
    wire N__48545;
    wire N__48540;
    wire N__48537;
    wire N__48534;
    wire N__48525;
    wire N__48524;
    wire N__48523;
    wire N__48520;
    wire N__48517;
    wire N__48514;
    wire N__48507;
    wire N__48504;
    wire N__48503;
    wire N__48502;
    wire N__48501;
    wire N__48498;
    wire N__48491;
    wire N__48486;
    wire N__48483;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48471;
    wire N__48468;
    wire N__48467;
    wire N__48464;
    wire N__48461;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48450;
    wire N__48447;
    wire N__48442;
    wire N__48439;
    wire N__48432;
    wire N__48429;
    wire N__48426;
    wire N__48425;
    wire N__48422;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48412;
    wire N__48405;
    wire N__48402;
    wire N__48399;
    wire N__48396;
    wire N__48393;
    wire N__48392;
    wire N__48389;
    wire N__48386;
    wire N__48385;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48373;
    wire N__48368;
    wire N__48365;
    wire N__48360;
    wire N__48357;
    wire N__48354;
    wire N__48353;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48336;
    wire N__48333;
    wire N__48330;
    wire N__48327;
    wire N__48324;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48314;
    wire N__48313;
    wire N__48310;
    wire N__48305;
    wire N__48304;
    wire N__48299;
    wire N__48296;
    wire N__48291;
    wire N__48288;
    wire N__48287;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48277;
    wire N__48270;
    wire N__48267;
    wire N__48264;
    wire N__48261;
    wire N__48258;
    wire N__48255;
    wire N__48254;
    wire N__48253;
    wire N__48252;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48244;
    wire N__48243;
    wire N__48242;
    wire N__48241;
    wire N__48240;
    wire N__48239;
    wire N__48238;
    wire N__48237;
    wire N__48236;
    wire N__48235;
    wire N__48234;
    wire N__48229;
    wire N__48228;
    wire N__48227;
    wire N__48226;
    wire N__48225;
    wire N__48224;
    wire N__48223;
    wire N__48222;
    wire N__48221;
    wire N__48220;
    wire N__48217;
    wire N__48216;
    wire N__48215;
    wire N__48214;
    wire N__48213;
    wire N__48212;
    wire N__48211;
    wire N__48210;
    wire N__48209;
    wire N__48208;
    wire N__48207;
    wire N__48206;
    wire N__48205;
    wire N__48202;
    wire N__48199;
    wire N__48198;
    wire N__48197;
    wire N__48196;
    wire N__48191;
    wire N__48188;
    wire N__48187;
    wire N__48186;
    wire N__48185;
    wire N__48184;
    wire N__48183;
    wire N__48182;
    wire N__48181;
    wire N__48180;
    wire N__48179;
    wire N__48170;
    wire N__48169;
    wire N__48168;
    wire N__48167;
    wire N__48166;
    wire N__48165;
    wire N__48164;
    wire N__48159;
    wire N__48154;
    wire N__48151;
    wire N__48142;
    wire N__48127;
    wire N__48110;
    wire N__48107;
    wire N__48104;
    wire N__48101;
    wire N__48098;
    wire N__48095;
    wire N__48094;
    wire N__48093;
    wire N__48092;
    wire N__48091;
    wire N__48088;
    wire N__48087;
    wire N__48086;
    wire N__48085;
    wire N__48084;
    wire N__48083;
    wire N__48082;
    wire N__48081;
    wire N__48080;
    wire N__48079;
    wire N__48074;
    wire N__48071;
    wire N__48068;
    wire N__48061;
    wire N__48056;
    wire N__48047;
    wire N__48044;
    wire N__48031;
    wire N__48016;
    wire N__48011;
    wire N__48010;
    wire N__48009;
    wire N__48008;
    wire N__48003;
    wire N__47998;
    wire N__47995;
    wire N__47990;
    wire N__47987;
    wire N__47984;
    wire N__47969;
    wire N__47956;
    wire N__47947;
    wire N__47940;
    wire N__47919;
    wire N__47918;
    wire N__47915;
    wire N__47912;
    wire N__47911;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47892;
    wire N__47889;
    wire N__47880;
    wire N__47879;
    wire N__47878;
    wire N__47877;
    wire N__47876;
    wire N__47875;
    wire N__47874;
    wire N__47873;
    wire N__47872;
    wire N__47871;
    wire N__47870;
    wire N__47867;
    wire N__47866;
    wire N__47865;
    wire N__47864;
    wire N__47863;
    wire N__47862;
    wire N__47861;
    wire N__47858;
    wire N__47857;
    wire N__47854;
    wire N__47853;
    wire N__47850;
    wire N__47849;
    wire N__47848;
    wire N__47847;
    wire N__47846;
    wire N__47843;
    wire N__47840;
    wire N__47839;
    wire N__47838;
    wire N__47837;
    wire N__47836;
    wire N__47835;
    wire N__47834;
    wire N__47831;
    wire N__47830;
    wire N__47827;
    wire N__47826;
    wire N__47823;
    wire N__47822;
    wire N__47821;
    wire N__47820;
    wire N__47819;
    wire N__47818;
    wire N__47817;
    wire N__47816;
    wire N__47815;
    wire N__47814;
    wire N__47813;
    wire N__47812;
    wire N__47811;
    wire N__47810;
    wire N__47809;
    wire N__47808;
    wire N__47807;
    wire N__47802;
    wire N__47801;
    wire N__47800;
    wire N__47799;
    wire N__47798;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47792;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47782;
    wire N__47769;
    wire N__47768;
    wire N__47763;
    wire N__47758;
    wire N__47757;
    wire N__47756;
    wire N__47755;
    wire N__47754;
    wire N__47751;
    wire N__47750;
    wire N__47747;
    wire N__47746;
    wire N__47745;
    wire N__47744;
    wire N__47743;
    wire N__47742;
    wire N__47741;
    wire N__47740;
    wire N__47739;
    wire N__47736;
    wire N__47733;
    wire N__47730;
    wire N__47729;
    wire N__47726;
    wire N__47725;
    wire N__47722;
    wire N__47721;
    wire N__47718;
    wire N__47701;
    wire N__47698;
    wire N__47697;
    wire N__47694;
    wire N__47693;
    wire N__47690;
    wire N__47689;
    wire N__47686;
    wire N__47685;
    wire N__47682;
    wire N__47681;
    wire N__47678;
    wire N__47677;
    wire N__47674;
    wire N__47673;
    wire N__47670;
    wire N__47669;
    wire N__47666;
    wire N__47665;
    wire N__47662;
    wire N__47661;
    wire N__47658;
    wire N__47657;
    wire N__47654;
    wire N__47653;
    wire N__47650;
    wire N__47649;
    wire N__47646;
    wire N__47645;
    wire N__47642;
    wire N__47641;
    wire N__47638;
    wire N__47631;
    wire N__47624;
    wire N__47623;
    wire N__47620;
    wire N__47619;
    wire N__47618;
    wire N__47617;
    wire N__47616;
    wire N__47615;
    wire N__47614;
    wire N__47613;
    wire N__47612;
    wire N__47611;
    wire N__47610;
    wire N__47607;
    wire N__47604;
    wire N__47597;
    wire N__47594;
    wire N__47591;
    wire N__47590;
    wire N__47589;
    wire N__47588;
    wire N__47587;
    wire N__47586;
    wire N__47585;
    wire N__47584;
    wire N__47579;
    wire N__47564;
    wire N__47547;
    wire N__47542;
    wire N__47527;
    wire N__47524;
    wire N__47507;
    wire N__47490;
    wire N__47473;
    wire N__47460;
    wire N__47455;
    wire N__47452;
    wire N__47445;
    wire N__47430;
    wire N__47429;
    wire N__47428;
    wire N__47427;
    wire N__47426;
    wire N__47423;
    wire N__47420;
    wire N__47419;
    wire N__47418;
    wire N__47407;
    wire N__47404;
    wire N__47403;
    wire N__47400;
    wire N__47399;
    wire N__47396;
    wire N__47395;
    wire N__47392;
    wire N__47391;
    wire N__47388;
    wire N__47387;
    wire N__47384;
    wire N__47383;
    wire N__47380;
    wire N__47379;
    wire N__47358;
    wire N__47355;
    wire N__47348;
    wire N__47335;
    wire N__47330;
    wire N__47327;
    wire N__47310;
    wire N__47297;
    wire N__47294;
    wire N__47277;
    wire N__47274;
    wire N__47273;
    wire N__47272;
    wire N__47269;
    wire N__47266;
    wire N__47263;
    wire N__47260;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47243;
    wire N__47240;
    wire N__47237;
    wire N__47234;
    wire N__47233;
    wire N__47232;
    wire N__47229;
    wire N__47226;
    wire N__47221;
    wire N__47218;
    wire N__47211;
    wire N__47208;
    wire N__47205;
    wire N__47202;
    wire N__47201;
    wire N__47198;
    wire N__47195;
    wire N__47190;
    wire N__47189;
    wire N__47184;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47174;
    wire N__47169;
    wire N__47166;
    wire N__47163;
    wire N__47162;
    wire N__47161;
    wire N__47160;
    wire N__47159;
    wire N__47158;
    wire N__47157;
    wire N__47156;
    wire N__47155;
    wire N__47154;
    wire N__47153;
    wire N__47152;
    wire N__47127;
    wire N__47124;
    wire N__47121;
    wire N__47120;
    wire N__47117;
    wire N__47114;
    wire N__47113;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47092;
    wire N__47089;
    wire N__47084;
    wire N__47081;
    wire N__47076;
    wire N__47075;
    wire N__47074;
    wire N__47071;
    wire N__47070;
    wire N__47069;
    wire N__47064;
    wire N__47061;
    wire N__47060;
    wire N__47059;
    wire N__47058;
    wire N__47057;
    wire N__47056;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47048;
    wire N__47047;
    wire N__47046;
    wire N__47045;
    wire N__47044;
    wire N__47043;
    wire N__47042;
    wire N__47041;
    wire N__47040;
    wire N__47039;
    wire N__47038;
    wire N__47037;
    wire N__47036;
    wire N__47035;
    wire N__47034;
    wire N__47033;
    wire N__47032;
    wire N__47031;
    wire N__47030;
    wire N__47029;
    wire N__47028;
    wire N__47027;
    wire N__47026;
    wire N__47025;
    wire N__47024;
    wire N__47023;
    wire N__47022;
    wire N__47021;
    wire N__47020;
    wire N__47017;
    wire N__47014;
    wire N__47007;
    wire N__47000;
    wire N__46995;
    wire N__46992;
    wire N__46991;
    wire N__46988;
    wire N__46979;
    wire N__46972;
    wire N__46971;
    wire N__46970;
    wire N__46969;
    wire N__46966;
    wire N__46965;
    wire N__46964;
    wire N__46961;
    wire N__46960;
    wire N__46959;
    wire N__46958;
    wire N__46957;
    wire N__46956;
    wire N__46955;
    wire N__46944;
    wire N__46943;
    wire N__46942;
    wire N__46941;
    wire N__46940;
    wire N__46937;
    wire N__46936;
    wire N__46935;
    wire N__46934;
    wire N__46933;
    wire N__46922;
    wire N__46921;
    wire N__46920;
    wire N__46919;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46913;
    wire N__46912;
    wire N__46903;
    wire N__46896;
    wire N__46889;
    wire N__46882;
    wire N__46881;
    wire N__46880;
    wire N__46879;
    wire N__46876;
    wire N__46875;
    wire N__46874;
    wire N__46867;
    wire N__46854;
    wire N__46853;
    wire N__46852;
    wire N__46851;
    wire N__46850;
    wire N__46849;
    wire N__46846;
    wire N__46835;
    wire N__46832;
    wire N__46831;
    wire N__46830;
    wire N__46827;
    wire N__46818;
    wire N__46817;
    wire N__46816;
    wire N__46815;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46808;
    wire N__46805;
    wire N__46798;
    wire N__46795;
    wire N__46782;
    wire N__46775;
    wire N__46772;
    wire N__46763;
    wire N__46760;
    wire N__46749;
    wire N__46744;
    wire N__46733;
    wire N__46728;
    wire N__46725;
    wire N__46724;
    wire N__46723;
    wire N__46722;
    wire N__46717;
    wire N__46712;
    wire N__46703;
    wire N__46696;
    wire N__46689;
    wire N__46686;
    wire N__46681;
    wire N__46676;
    wire N__46671;
    wire N__46664;
    wire N__46661;
    wire N__46658;
    wire N__46653;
    wire N__46648;
    wire N__46639;
    wire N__46634;
    wire N__46629;
    wire N__46626;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46604;
    wire N__46601;
    wire N__46598;
    wire N__46595;
    wire N__46590;
    wire N__46587;
    wire N__46584;
    wire N__46581;
    wire N__46578;
    wire N__46577;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46557;
    wire N__46554;
    wire N__46553;
    wire N__46550;
    wire N__46547;
    wire N__46544;
    wire N__46539;
    wire N__46536;
    wire N__46533;
    wire N__46530;
    wire N__46529;
    wire N__46526;
    wire N__46525;
    wire N__46522;
    wire N__46519;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46507;
    wire N__46504;
    wire N__46499;
    wire N__46494;
    wire N__46491;
    wire N__46490;
    wire N__46487;
    wire N__46484;
    wire N__46483;
    wire N__46480;
    wire N__46477;
    wire N__46474;
    wire N__46469;
    wire N__46464;
    wire N__46461;
    wire N__46460;
    wire N__46459;
    wire N__46458;
    wire N__46455;
    wire N__46452;
    wire N__46447;
    wire N__46440;
    wire N__46439;
    wire N__46436;
    wire N__46433;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46418;
    wire N__46413;
    wire N__46412;
    wire N__46411;
    wire N__46410;
    wire N__46409;
    wire N__46408;
    wire N__46407;
    wire N__46406;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46377;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46359;
    wire N__46354;
    wire N__46351;
    wire N__46348;
    wire N__46343;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46322;
    wire N__46319;
    wire N__46316;
    wire N__46315;
    wire N__46310;
    wire N__46307;
    wire N__46304;
    wire N__46299;
    wire N__46296;
    wire N__46293;
    wire N__46292;
    wire N__46289;
    wire N__46286;
    wire N__46285;
    wire N__46280;
    wire N__46277;
    wire N__46274;
    wire N__46269;
    wire N__46266;
    wire N__46265;
    wire N__46260;
    wire N__46259;
    wire N__46256;
    wire N__46253;
    wire N__46250;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46238;
    wire N__46237;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46217;
    wire N__46214;
    wire N__46209;
    wire N__46206;
    wire N__46205;
    wire N__46202;
    wire N__46199;
    wire N__46196;
    wire N__46193;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46170;
    wire N__46167;
    wire N__46166;
    wire N__46161;
    wire N__46160;
    wire N__46157;
    wire N__46154;
    wire N__46151;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46139;
    wire N__46136;
    wire N__46133;
    wire N__46132;
    wire N__46127;
    wire N__46124;
    wire N__46121;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46106;
    wire N__46103;
    wire N__46100;
    wire N__46097;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46085;
    wire N__46082;
    wire N__46079;
    wire N__46078;
    wire N__46073;
    wire N__46070;
    wire N__46067;
    wire N__46062;
    wire N__46059;
    wire N__46058;
    wire N__46055;
    wire N__46052;
    wire N__46047;
    wire N__46046;
    wire N__46043;
    wire N__46040;
    wire N__46037;
    wire N__46032;
    wire N__46029;
    wire N__46026;
    wire N__46025;
    wire N__46022;
    wire N__46019;
    wire N__46018;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__46002;
    wire N__45999;
    wire N__45998;
    wire N__45997;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45972;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45964;
    wire N__45961;
    wire N__45958;
    wire N__45955;
    wire N__45952;
    wire N__45949;
    wire N__45942;
    wire N__45939;
    wire N__45938;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45926;
    wire N__45925;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45902;
    wire N__45899;
    wire N__45896;
    wire N__45895;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45879;
    wire N__45876;
    wire N__45873;
    wire N__45872;
    wire N__45869;
    wire N__45866;
    wire N__45865;
    wire N__45860;
    wire N__45857;
    wire N__45854;
    wire N__45849;
    wire N__45846;
    wire N__45843;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45835;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45819;
    wire N__45816;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45804;
    wire N__45803;
    wire N__45800;
    wire N__45797;
    wire N__45794;
    wire N__45789;
    wire N__45786;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45774;
    wire N__45773;
    wire N__45770;
    wire N__45767;
    wire N__45764;
    wire N__45759;
    wire N__45756;
    wire N__45755;
    wire N__45750;
    wire N__45749;
    wire N__45746;
    wire N__45743;
    wire N__45740;
    wire N__45735;
    wire N__45732;
    wire N__45731;
    wire N__45726;
    wire N__45725;
    wire N__45722;
    wire N__45719;
    wire N__45716;
    wire N__45711;
    wire N__45708;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45694;
    wire N__45691;
    wire N__45688;
    wire N__45685;
    wire N__45682;
    wire N__45679;
    wire N__45672;
    wire N__45669;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45656;
    wire N__45655;
    wire N__45652;
    wire N__45649;
    wire N__45646;
    wire N__45643;
    wire N__45640;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45619;
    wire N__45614;
    wire N__45611;
    wire N__45608;
    wire N__45603;
    wire N__45600;
    wire N__45599;
    wire N__45594;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45579;
    wire N__45576;
    wire N__45575;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45563;
    wire N__45562;
    wire N__45559;
    wire N__45556;
    wire N__45551;
    wire N__45546;
    wire N__45545;
    wire N__45544;
    wire N__45541;
    wire N__45536;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45515;
    wire N__45514;
    wire N__45511;
    wire N__45508;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45481;
    wire N__45474;
    wire N__45471;
    wire N__45468;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45456;
    wire N__45455;
    wire N__45452;
    wire N__45447;
    wire N__45444;
    wire N__45443;
    wire N__45442;
    wire N__45441;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45414;
    wire N__45411;
    wire N__45408;
    wire N__45407;
    wire N__45404;
    wire N__45401;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45376;
    wire N__45373;
    wire N__45370;
    wire N__45367;
    wire N__45364;
    wire N__45361;
    wire N__45354;
    wire N__45353;
    wire N__45352;
    wire N__45349;
    wire N__45346;
    wire N__45343;
    wire N__45342;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45328;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45295;
    wire N__45292;
    wire N__45289;
    wire N__45286;
    wire N__45281;
    wire N__45276;
    wire N__45273;
    wire N__45272;
    wire N__45267;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45252;
    wire N__45249;
    wire N__45248;
    wire N__45243;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45233;
    wire N__45228;
    wire N__45225;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45212;
    wire N__45209;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45192;
    wire N__45191;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45178;
    wire N__45173;
    wire N__45172;
    wire N__45167;
    wire N__45164;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45146;
    wire N__45143;
    wire N__45140;
    wire N__45139;
    wire N__45136;
    wire N__45133;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45095;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45083;
    wire N__45082;
    wire N__45079;
    wire N__45076;
    wire N__45071;
    wire N__45066;
    wire N__45065;
    wire N__45064;
    wire N__45061;
    wire N__45056;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45038;
    wire N__45035;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45020;
    wire N__45015;
    wire N__45014;
    wire N__45013;
    wire N__45010;
    wire N__45007;
    wire N__45004;
    wire N__45003;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44980;
    wire N__44973;
    wire N__44972;
    wire N__44969;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44955;
    wire N__44952;
    wire N__44949;
    wire N__44948;
    wire N__44947;
    wire N__44944;
    wire N__44941;
    wire N__44938;
    wire N__44935;
    wire N__44928;
    wire N__44927;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44915;
    wire N__44914;
    wire N__44911;
    wire N__44908;
    wire N__44905;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44873;
    wire N__44872;
    wire N__44871;
    wire N__44870;
    wire N__44869;
    wire N__44868;
    wire N__44867;
    wire N__44866;
    wire N__44865;
    wire N__44864;
    wire N__44863;
    wire N__44854;
    wire N__44853;
    wire N__44852;
    wire N__44851;
    wire N__44850;
    wire N__44849;
    wire N__44848;
    wire N__44847;
    wire N__44846;
    wire N__44837;
    wire N__44828;
    wire N__44827;
    wire N__44826;
    wire N__44825;
    wire N__44824;
    wire N__44823;
    wire N__44822;
    wire N__44821;
    wire N__44820;
    wire N__44819;
    wire N__44818;
    wire N__44815;
    wire N__44806;
    wire N__44797;
    wire N__44792;
    wire N__44787;
    wire N__44778;
    wire N__44769;
    wire N__44762;
    wire N__44755;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44739;
    wire N__44736;
    wire N__44733;
    wire N__44730;
    wire N__44729;
    wire N__44726;
    wire N__44723;
    wire N__44720;
    wire N__44715;
    wire N__44714;
    wire N__44713;
    wire N__44710;
    wire N__44707;
    wire N__44706;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44694;
    wire N__44691;
    wire N__44686;
    wire N__44683;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44667;
    wire N__44664;
    wire N__44663;
    wire N__44662;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44636;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44624;
    wire N__44621;
    wire N__44618;
    wire N__44613;
    wire N__44612;
    wire N__44611;
    wire N__44608;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44589;
    wire N__44588;
    wire N__44585;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44574;
    wire N__44571;
    wire N__44566;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44554;
    wire N__44547;
    wire N__44546;
    wire N__44545;
    wire N__44542;
    wire N__44537;
    wire N__44534;
    wire N__44531;
    wire N__44530;
    wire N__44525;
    wire N__44522;
    wire N__44517;
    wire N__44514;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44502;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44490;
    wire N__44487;
    wire N__44484;
    wire N__44481;
    wire N__44478;
    wire N__44477;
    wire N__44476;
    wire N__44473;
    wire N__44470;
    wire N__44465;
    wire N__44460;
    wire N__44459;
    wire N__44458;
    wire N__44455;
    wire N__44452;
    wire N__44447;
    wire N__44442;
    wire N__44441;
    wire N__44436;
    wire N__44433;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44421;
    wire N__44418;
    wire N__44417;
    wire N__44416;
    wire N__44413;
    wire N__44408;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44398;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44364;
    wire N__44363;
    wire N__44358;
    wire N__44355;
    wire N__44354;
    wire N__44351;
    wire N__44348;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44332;
    wire N__44325;
    wire N__44322;
    wire N__44321;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44310;
    wire N__44307;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44289;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44277;
    wire N__44276;
    wire N__44273;
    wire N__44270;
    wire N__44267;
    wire N__44262;
    wire N__44259;
    wire N__44258;
    wire N__44255;
    wire N__44252;
    wire N__44247;
    wire N__44246;
    wire N__44243;
    wire N__44240;
    wire N__44237;
    wire N__44232;
    wire N__44229;
    wire N__44228;
    wire N__44223;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44201;
    wire N__44198;
    wire N__44195;
    wire N__44194;
    wire N__44189;
    wire N__44186;
    wire N__44183;
    wire N__44178;
    wire N__44175;
    wire N__44174;
    wire N__44171;
    wire N__44168;
    wire N__44165;
    wire N__44162;
    wire N__44161;
    wire N__44156;
    wire N__44153;
    wire N__44150;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44138;
    wire N__44135;
    wire N__44132;
    wire N__44131;
    wire N__44128;
    wire N__44125;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44109;
    wire N__44106;
    wire N__44103;
    wire N__44102;
    wire N__44099;
    wire N__44096;
    wire N__44095;
    wire N__44090;
    wire N__44087;
    wire N__44084;
    wire N__44079;
    wire N__44076;
    wire N__44075;
    wire N__44070;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44048;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44034;
    wire N__44033;
    wire N__44028;
    wire N__44027;
    wire N__44024;
    wire N__44021;
    wire N__44018;
    wire N__44013;
    wire N__44010;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__43998;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43983;
    wire N__43980;
    wire N__43979;
    wire N__43976;
    wire N__43973;
    wire N__43968;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43958;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43939;
    wire N__43934;
    wire N__43931;
    wire N__43928;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43909;
    wire N__43904;
    wire N__43901;
    wire N__43898;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43886;
    wire N__43883;
    wire N__43880;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43857;
    wire N__43854;
    wire N__43853;
    wire N__43848;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43833;
    wire N__43830;
    wire N__43829;
    wire N__43824;
    wire N__43823;
    wire N__43820;
    wire N__43817;
    wire N__43814;
    wire N__43809;
    wire N__43806;
    wire N__43805;
    wire N__43802;
    wire N__43799;
    wire N__43794;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43779;
    wire N__43776;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43764;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43754;
    wire N__43749;
    wire N__43746;
    wire N__43743;
    wire N__43742;
    wire N__43739;
    wire N__43736;
    wire N__43735;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43719;
    wire N__43716;
    wire N__43715;
    wire N__43710;
    wire N__43709;
    wire N__43706;
    wire N__43703;
    wire N__43700;
    wire N__43695;
    wire N__43692;
    wire N__43691;
    wire N__43686;
    wire N__43685;
    wire N__43682;
    wire N__43679;
    wire N__43676;
    wire N__43671;
    wire N__43668;
    wire N__43667;
    wire N__43664;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43654;
    wire N__43649;
    wire N__43646;
    wire N__43643;
    wire N__43638;
    wire N__43635;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43618;
    wire N__43615;
    wire N__43612;
    wire N__43609;
    wire N__43604;
    wire N__43599;
    wire N__43596;
    wire N__43593;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43585;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43569;
    wire N__43566;
    wire N__43565;
    wire N__43560;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43519;
    wire N__43514;
    wire N__43511;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43501;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43485;
    wire N__43484;
    wire N__43481;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43471;
    wire N__43470;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43452;
    wire N__43449;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43383;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43375;
    wire N__43372;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43354;
    wire N__43349;
    wire N__43344;
    wire N__43343;
    wire N__43340;
    wire N__43337;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43319;
    wire N__43314;
    wire N__43311;
    wire N__43308;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43298;
    wire N__43295;
    wire N__43292;
    wire N__43289;
    wire N__43288;
    wire N__43283;
    wire N__43280;
    wire N__43277;
    wire N__43272;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43256;
    wire N__43253;
    wire N__43250;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43240;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43205;
    wire N__43202;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43191;
    wire N__43188;
    wire N__43183;
    wire N__43180;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43140;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43103;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43092;
    wire N__43089;
    wire N__43084;
    wire N__43081;
    wire N__43074;
    wire N__43071;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43061;
    wire N__43058;
    wire N__43055;
    wire N__43052;
    wire N__43049;
    wire N__43048;
    wire N__43043;
    wire N__43040;
    wire N__43039;
    wire N__43036;
    wire N__43033;
    wire N__43030;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42987;
    wire N__42984;
    wire N__42979;
    wire N__42976;
    wire N__42969;
    wire N__42966;
    wire N__42963;
    wire N__42960;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42940;
    wire N__42939;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42897;
    wire N__42896;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42879;
    wire N__42876;
    wire N__42873;
    wire N__42870;
    wire N__42867;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42845;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42818;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42808;
    wire N__42805;
    wire N__42800;
    wire N__42799;
    wire N__42794;
    wire N__42791;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42777;
    wire N__42774;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42759;
    wire N__42758;
    wire N__42757;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42738;
    wire N__42731;
    wire N__42728;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42714;
    wire N__42713;
    wire N__42710;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42698;
    wire N__42697;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42687;
    wire N__42684;
    wire N__42679;
    wire N__42676;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42641;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42631;
    wire N__42628;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42605;
    wire N__42602;
    wire N__42599;
    wire N__42598;
    wire N__42593;
    wire N__42590;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42580;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42551;
    wire N__42550;
    wire N__42547;
    wire N__42544;
    wire N__42541;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42515;
    wire N__42512;
    wire N__42509;
    wire N__42508;
    wire N__42505;
    wire N__42502;
    wire N__42499;
    wire N__42492;
    wire N__42489;
    wire N__42486;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42478;
    wire N__42473;
    wire N__42470;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42458;
    wire N__42457;
    wire N__42454;
    wire N__42451;
    wire N__42448;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42431;
    wire N__42428;
    wire N__42423;
    wire N__42420;
    wire N__42419;
    wire N__42418;
    wire N__42415;
    wire N__42412;
    wire N__42409;
    wire N__42406;
    wire N__42401;
    wire N__42398;
    wire N__42393;
    wire N__42390;
    wire N__42389;
    wire N__42388;
    wire N__42385;
    wire N__42382;
    wire N__42379;
    wire N__42376;
    wire N__42373;
    wire N__42370;
    wire N__42367;
    wire N__42362;
    wire N__42357;
    wire N__42354;
    wire N__42353;
    wire N__42352;
    wire N__42349;
    wire N__42346;
    wire N__42343;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42314;
    wire N__42311;
    wire N__42310;
    wire N__42307;
    wire N__42304;
    wire N__42301;
    wire N__42298;
    wire N__42295;
    wire N__42292;
    wire N__42289;
    wire N__42282;
    wire N__42279;
    wire N__42278;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42268;
    wire N__42265;
    wire N__42262;
    wire N__42259;
    wire N__42252;
    wire N__42249;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42236;
    wire N__42235;
    wire N__42230;
    wire N__42227;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42212;
    wire N__42211;
    wire N__42208;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42196;
    wire N__42193;
    wire N__42188;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42176;
    wire N__42175;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42157;
    wire N__42152;
    wire N__42149;
    wire N__42144;
    wire N__42141;
    wire N__42140;
    wire N__42137;
    wire N__42136;
    wire N__42133;
    wire N__42130;
    wire N__42127;
    wire N__42124;
    wire N__42121;
    wire N__42118;
    wire N__42113;
    wire N__42110;
    wire N__42105;
    wire N__42102;
    wire N__42099;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42089;
    wire N__42086;
    wire N__42085;
    wire N__42082;
    wire N__42079;
    wire N__42076;
    wire N__42073;
    wire N__42068;
    wire N__42065;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42053;
    wire N__42050;
    wire N__42047;
    wire N__42044;
    wire N__42041;
    wire N__42040;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42024;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42008;
    wire N__42005;
    wire N__42002;
    wire N__41999;
    wire N__41996;
    wire N__41995;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41972;
    wire N__41969;
    wire N__41966;
    wire N__41965;
    wire N__41960;
    wire N__41957;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41936;
    wire N__41935;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41882;
    wire N__41879;
    wire N__41876;
    wire N__41873;
    wire N__41870;
    wire N__41867;
    wire N__41864;
    wire N__41861;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41841;
    wire N__41838;
    wire N__41837;
    wire N__41836;
    wire N__41833;
    wire N__41828;
    wire N__41827;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41809;
    wire N__41802;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41767;
    wire N__41762;
    wire N__41759;
    wire N__41754;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41744;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41727;
    wire N__41724;
    wire N__41721;
    wire N__41718;
    wire N__41717;
    wire N__41716;
    wire N__41713;
    wire N__41708;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41696;
    wire N__41695;
    wire N__41692;
    wire N__41687;
    wire N__41682;
    wire N__41679;
    wire N__41678;
    wire N__41677;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41665;
    wire N__41662;
    wire N__41655;
    wire N__41652;
    wire N__41651;
    wire N__41648;
    wire N__41645;
    wire N__41640;
    wire N__41639;
    wire N__41634;
    wire N__41631;
    wire N__41630;
    wire N__41625;
    wire N__41624;
    wire N__41623;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41609;
    wire N__41604;
    wire N__41601;
    wire N__41598;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41586;
    wire N__41585;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41575;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41559;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41551;
    wire N__41550;
    wire N__41547;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41533;
    wire N__41526;
    wire N__41525;
    wire N__41522;
    wire N__41519;
    wire N__41514;
    wire N__41513;
    wire N__41510;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41475;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41461;
    wire N__41456;
    wire N__41453;
    wire N__41450;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41433;
    wire N__41432;
    wire N__41431;
    wire N__41430;
    wire N__41427;
    wire N__41424;
    wire N__41421;
    wire N__41418;
    wire N__41413;
    wire N__41408;
    wire N__41405;
    wire N__41400;
    wire N__41397;
    wire N__41396;
    wire N__41395;
    wire N__41392;
    wire N__41389;
    wire N__41386;
    wire N__41383;
    wire N__41376;
    wire N__41375;
    wire N__41374;
    wire N__41371;
    wire N__41368;
    wire N__41367;
    wire N__41364;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41343;
    wire N__41342;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41319;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41294;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41279;
    wire N__41278;
    wire N__41277;
    wire N__41276;
    wire N__41275;
    wire N__41274;
    wire N__41273;
    wire N__41272;
    wire N__41271;
    wire N__41270;
    wire N__41269;
    wire N__41266;
    wire N__41265;
    wire N__41264;
    wire N__41263;
    wire N__41254;
    wire N__41253;
    wire N__41252;
    wire N__41251;
    wire N__41250;
    wire N__41249;
    wire N__41248;
    wire N__41247;
    wire N__41246;
    wire N__41245;
    wire N__41244;
    wire N__41243;
    wire N__41242;
    wire N__41235;
    wire N__41226;
    wire N__41223;
    wire N__41216;
    wire N__41215;
    wire N__41214;
    wire N__41213;
    wire N__41212;
    wire N__41211;
    wire N__41208;
    wire N__41199;
    wire N__41190;
    wire N__41181;
    wire N__41178;
    wire N__41175;
    wire N__41172;
    wire N__41169;
    wire N__41166;
    wire N__41157;
    wire N__41144;
    wire N__41141;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41120;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41081;
    wire N__41078;
    wire N__41077;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41061;
    wire N__41058;
    wire N__41057;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41042;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41024;
    wire N__41023;
    wire N__41020;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41001;
    wire N__40998;
    wire N__40997;
    wire N__40996;
    wire N__40993;
    wire N__40988;
    wire N__40987;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40961;
    wire N__40960;
    wire N__40957;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40947;
    wire N__40940;
    wire N__40937;
    wire N__40934;
    wire N__40929;
    wire N__40926;
    wire N__40925;
    wire N__40922;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40890;
    wire N__40887;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40866;
    wire N__40863;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40847;
    wire N__40846;
    wire N__40841;
    wire N__40838;
    wire N__40835;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40823;
    wire N__40822;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40806;
    wire N__40803;
    wire N__40802;
    wire N__40799;
    wire N__40796;
    wire N__40791;
    wire N__40788;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40776;
    wire N__40773;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40761;
    wire N__40758;
    wire N__40757;
    wire N__40754;
    wire N__40751;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40734;
    wire N__40733;
    wire N__40728;
    wire N__40727;
    wire N__40724;
    wire N__40721;
    wire N__40718;
    wire N__40713;
    wire N__40710;
    wire N__40709;
    wire N__40704;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40682;
    wire N__40679;
    wire N__40676;
    wire N__40671;
    wire N__40668;
    wire N__40667;
    wire N__40664;
    wire N__40661;
    wire N__40656;
    wire N__40653;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40641;
    wire N__40638;
    wire N__40637;
    wire N__40634;
    wire N__40631;
    wire N__40626;
    wire N__40623;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40611;
    wire N__40608;
    wire N__40607;
    wire N__40604;
    wire N__40601;
    wire N__40596;
    wire N__40593;
    wire N__40592;
    wire N__40589;
    wire N__40586;
    wire N__40581;
    wire N__40578;
    wire N__40577;
    wire N__40574;
    wire N__40571;
    wire N__40566;
    wire N__40563;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40552;
    wire N__40549;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40525;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40478;
    wire N__40477;
    wire N__40474;
    wire N__40469;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40440;
    wire N__40437;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40418;
    wire N__40415;
    wire N__40414;
    wire N__40411;
    wire N__40408;
    wire N__40405;
    wire N__40398;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40325;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40317;
    wire N__40314;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40298;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40249;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40237;
    wire N__40234;
    wire N__40229;
    wire N__40224;
    wire N__40221;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40204;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40159;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40147;
    wire N__40142;
    wire N__40139;
    wire N__40134;
    wire N__40131;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40095;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40085;
    wire N__40082;
    wire N__40081;
    wire N__40080;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40037;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40008;
    wire N__40005;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39759;
    wire N__39756;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39720;
    wire N__39717;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39695;
    wire N__39694;
    wire N__39693;
    wire N__39690;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39657;
    wire N__39654;
    wire N__39653;
    wire N__39650;
    wire N__39649;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39633;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39615;
    wire N__39612;
    wire N__39611;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39600;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39584;
    wire N__39581;
    wire N__39578;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39564;
    wire N__39563;
    wire N__39562;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39550;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39534;
    wire N__39533;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39525;
    wire N__39522;
    wire N__39517;
    wire N__39512;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39464;
    wire N__39461;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39450;
    wire N__39447;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39396;
    wire N__39393;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39371;
    wire N__39370;
    wire N__39365;
    wire N__39362;
    wire N__39357;
    wire N__39354;
    wire N__39353;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39338;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39321;
    wire N__39318;
    wire N__39317;
    wire N__39316;
    wire N__39315;
    wire N__39310;
    wire N__39307;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39289;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39272;
    wire N__39269;
    wire N__39268;
    wire N__39265;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39247;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39066;
    wire N__39063;
    wire N__39062;
    wire N__39061;
    wire N__39060;
    wire N__39059;
    wire N__39052;
    wire N__39047;
    wire N__39044;
    wire N__39039;
    wire N__39036;
    wire N__39035;
    wire N__39030;
    wire N__39027;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39019;
    wire N__39018;
    wire N__39013;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38985;
    wire N__38984;
    wire N__38981;
    wire N__38980;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38907;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38861;
    wire N__38860;
    wire N__38859;
    wire N__38858;
    wire N__38857;
    wire N__38856;
    wire N__38855;
    wire N__38854;
    wire N__38853;
    wire N__38852;
    wire N__38851;
    wire N__38850;
    wire N__38849;
    wire N__38848;
    wire N__38845;
    wire N__38838;
    wire N__38829;
    wire N__38828;
    wire N__38825;
    wire N__38824;
    wire N__38821;
    wire N__38820;
    wire N__38817;
    wire N__38816;
    wire N__38815;
    wire N__38812;
    wire N__38811;
    wire N__38808;
    wire N__38807;
    wire N__38804;
    wire N__38803;
    wire N__38800;
    wire N__38793;
    wire N__38778;
    wire N__38763;
    wire N__38762;
    wire N__38761;
    wire N__38760;
    wire N__38759;
    wire N__38758;
    wire N__38757;
    wire N__38756;
    wire N__38755;
    wire N__38754;
    wire N__38753;
    wire N__38750;
    wire N__38749;
    wire N__38748;
    wire N__38747;
    wire N__38746;
    wire N__38743;
    wire N__38740;
    wire N__38737;
    wire N__38736;
    wire N__38733;
    wire N__38732;
    wire N__38729;
    wire N__38728;
    wire N__38725;
    wire N__38724;
    wire N__38721;
    wire N__38718;
    wire N__38713;
    wire N__38710;
    wire N__38709;
    wire N__38708;
    wire N__38707;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38693;
    wire N__38690;
    wire N__38689;
    wire N__38686;
    wire N__38685;
    wire N__38682;
    wire N__38681;
    wire N__38680;
    wire N__38679;
    wire N__38678;
    wire N__38677;
    wire N__38676;
    wire N__38675;
    wire N__38674;
    wire N__38673;
    wire N__38672;
    wire N__38671;
    wire N__38670;
    wire N__38667;
    wire N__38662;
    wire N__38645;
    wire N__38638;
    wire N__38635;
    wire N__38630;
    wire N__38627;
    wire N__38622;
    wire N__38619;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38583;
    wire N__38574;
    wire N__38573;
    wire N__38572;
    wire N__38565;
    wire N__38556;
    wire N__38553;
    wire N__38548;
    wire N__38535;
    wire N__38532;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38516;
    wire N__38509;
    wire N__38502;
    wire N__38499;
    wire N__38498;
    wire N__38497;
    wire N__38496;
    wire N__38495;
    wire N__38494;
    wire N__38493;
    wire N__38492;
    wire N__38491;
    wire N__38490;
    wire N__38489;
    wire N__38486;
    wire N__38485;
    wire N__38480;
    wire N__38479;
    wire N__38476;
    wire N__38471;
    wire N__38468;
    wire N__38467;
    wire N__38464;
    wire N__38463;
    wire N__38462;
    wire N__38461;
    wire N__38460;
    wire N__38459;
    wire N__38458;
    wire N__38457;
    wire N__38456;
    wire N__38455;
    wire N__38454;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38432;
    wire N__38431;
    wire N__38430;
    wire N__38429;
    wire N__38428;
    wire N__38427;
    wire N__38426;
    wire N__38419;
    wire N__38406;
    wire N__38393;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38374;
    wire N__38365;
    wire N__38358;
    wire N__38349;
    wire N__38340;
    wire N__38335;
    wire N__38332;
    wire N__38327;
    wire N__38322;
    wire N__38321;
    wire N__38320;
    wire N__38317;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38297;
    wire N__38292;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38280;
    wire N__38277;
    wire N__38276;
    wire N__38273;
    wire N__38272;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38253;
    wire N__38250;
    wire N__38249;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38208;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38196;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38142;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37902;
    wire N__37901;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37886;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37857;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37758;
    wire N__37757;
    wire N__37754;
    wire N__37753;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37737;
    wire N__37736;
    wire N__37733;
    wire N__37732;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37703;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37691;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37679;
    wire N__37676;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37659;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37643;
    wire N__37642;
    wire N__37641;
    wire N__37640;
    wire N__37639;
    wire N__37638;
    wire N__37635;
    wire N__37634;
    wire N__37631;
    wire N__37630;
    wire N__37629;
    wire N__37628;
    wire N__37627;
    wire N__37626;
    wire N__37625;
    wire N__37624;
    wire N__37623;
    wire N__37622;
    wire N__37621;
    wire N__37620;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37612;
    wire N__37611;
    wire N__37610;
    wire N__37609;
    wire N__37608;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37590;
    wire N__37589;
    wire N__37588;
    wire N__37587;
    wire N__37586;
    wire N__37585;
    wire N__37584;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37568;
    wire N__37559;
    wire N__37558;
    wire N__37557;
    wire N__37556;
    wire N__37555;
    wire N__37548;
    wire N__37543;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37520;
    wire N__37519;
    wire N__37518;
    wire N__37515;
    wire N__37510;
    wire N__37509;
    wire N__37508;
    wire N__37507;
    wire N__37506;
    wire N__37503;
    wire N__37496;
    wire N__37487;
    wire N__37478;
    wire N__37469;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37430;
    wire N__37427;
    wire N__37416;
    wire N__37409;
    wire N__37404;
    wire N__37397;
    wire N__37392;
    wire N__37389;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37337;
    wire N__37332;
    wire N__37329;
    wire N__37328;
    wire N__37327;
    wire N__37324;
    wire N__37319;
    wire N__37314;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37302;
    wire N__37299;
    wire N__37298;
    wire N__37297;
    wire N__37294;
    wire N__37289;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37262;
    wire N__37259;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37242;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37221;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37200;
    wire N__37199;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37184;
    wire N__37179;
    wire N__37178;
    wire N__37177;
    wire N__37174;
    wire N__37169;
    wire N__37164;
    wire N__37163;
    wire N__37160;
    wire N__37159;
    wire N__37156;
    wire N__37151;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37130;
    wire N__37127;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37115;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37098;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37067;
    wire N__37064;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37052;
    wire N__37047;
    wire N__37044;
    wire N__37041;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37029;
    wire N__37026;
    wire N__37023;
    wire N__37020;
    wire N__37017;
    wire N__37014;
    wire N__37013;
    wire N__37012;
    wire N__37011;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__36997;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36981;
    wire N__36980;
    wire N__36979;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36954;
    wire N__36953;
    wire N__36950;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36911;
    wire N__36910;
    wire N__36907;
    wire N__36902;
    wire N__36897;
    wire N__36894;
    wire N__36893;
    wire N__36888;
    wire N__36885;
    wire N__36882;
    wire N__36881;
    wire N__36880;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36852;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36774;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36763;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36733;
    wire N__36728;
    wire N__36723;
    wire N__36722;
    wire N__36721;
    wire N__36720;
    wire N__36719;
    wire N__36718;
    wire N__36715;
    wire N__36714;
    wire N__36713;
    wire N__36712;
    wire N__36711;
    wire N__36708;
    wire N__36705;
    wire N__36704;
    wire N__36703;
    wire N__36702;
    wire N__36701;
    wire N__36700;
    wire N__36695;
    wire N__36692;
    wire N__36691;
    wire N__36690;
    wire N__36689;
    wire N__36688;
    wire N__36687;
    wire N__36686;
    wire N__36683;
    wire N__36682;
    wire N__36681;
    wire N__36680;
    wire N__36679;
    wire N__36678;
    wire N__36677;
    wire N__36676;
    wire N__36675;
    wire N__36674;
    wire N__36673;
    wire N__36672;
    wire N__36671;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36659;
    wire N__36652;
    wire N__36651;
    wire N__36650;
    wire N__36649;
    wire N__36646;
    wire N__36645;
    wire N__36642;
    wire N__36641;
    wire N__36640;
    wire N__36639;
    wire N__36638;
    wire N__36637;
    wire N__36636;
    wire N__36635;
    wire N__36634;
    wire N__36633;
    wire N__36632;
    wire N__36631;
    wire N__36630;
    wire N__36625;
    wire N__36620;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36603;
    wire N__36602;
    wire N__36599;
    wire N__36598;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36586;
    wire N__36573;
    wire N__36570;
    wire N__36565;
    wire N__36562;
    wire N__36561;
    wire N__36560;
    wire N__36559;
    wire N__36558;
    wire N__36557;
    wire N__36556;
    wire N__36555;
    wire N__36550;
    wire N__36547;
    wire N__36546;
    wire N__36545;
    wire N__36544;
    wire N__36543;
    wire N__36542;
    wire N__36539;
    wire N__36530;
    wire N__36527;
    wire N__36518;
    wire N__36513;
    wire N__36506;
    wire N__36503;
    wire N__36498;
    wire N__36491;
    wire N__36484;
    wire N__36479;
    wire N__36478;
    wire N__36477;
    wire N__36474;
    wire N__36473;
    wire N__36472;
    wire N__36471;
    wire N__36470;
    wire N__36469;
    wire N__36468;
    wire N__36467;
    wire N__36466;
    wire N__36465;
    wire N__36464;
    wire N__36463;
    wire N__36462;
    wire N__36457;
    wire N__36454;
    wire N__36451;
    wire N__36446;
    wire N__36439;
    wire N__36432;
    wire N__36423;
    wire N__36418;
    wire N__36417;
    wire N__36416;
    wire N__36415;
    wire N__36414;
    wire N__36413;
    wire N__36412;
    wire N__36411;
    wire N__36410;
    wire N__36409;
    wire N__36408;
    wire N__36407;
    wire N__36406;
    wire N__36401;
    wire N__36394;
    wire N__36391;
    wire N__36378;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36346;
    wire N__36341;
    wire N__36330;
    wire N__36327;
    wire N__36318;
    wire N__36311;
    wire N__36302;
    wire N__36291;
    wire N__36284;
    wire N__36273;
    wire N__36264;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36209;
    wire N__36204;
    wire N__36201;
    wire N__36198;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36192;
    wire N__36189;
    wire N__36184;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36159;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36147;
    wire N__36144;
    wire N__36141;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36048;
    wire N__36045;
    wire N__36042;
    wire N__36039;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35805;
    wire N__35802;
    wire N__35799;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35784;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35730;
    wire N__35727;
    wire N__35724;
    wire N__35721;
    wire N__35718;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35710;
    wire N__35707;
    wire N__35706;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35691;
    wire N__35688;
    wire N__35679;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35664;
    wire N__35661;
    wire N__35660;
    wire N__35657;
    wire N__35656;
    wire N__35655;
    wire N__35652;
    wire N__35649;
    wire N__35646;
    wire N__35643;
    wire N__35638;
    wire N__35635;
    wire N__35632;
    wire N__35629;
    wire N__35622;
    wire N__35621;
    wire N__35620;
    wire N__35619;
    wire N__35618;
    wire N__35613;
    wire N__35606;
    wire N__35603;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35582;
    wire N__35581;
    wire N__35578;
    wire N__35575;
    wire N__35570;
    wire N__35565;
    wire N__35562;
    wire N__35561;
    wire N__35560;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35544;
    wire N__35541;
    wire N__35540;
    wire N__35539;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35523;
    wire N__35520;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35484;
    wire N__35481;
    wire N__35478;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35400;
    wire N__35397;
    wire N__35396;
    wire N__35395;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35379;
    wire N__35376;
    wire N__35375;
    wire N__35372;
    wire N__35371;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35355;
    wire N__35352;
    wire N__35351;
    wire N__35350;
    wire N__35347;
    wire N__35342;
    wire N__35337;
    wire N__35334;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35322;
    wire N__35319;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35307;
    wire N__35304;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35292;
    wire N__35289;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35277;
    wire N__35274;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35262;
    wire N__35259;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35223;
    wire N__35220;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35199;
    wire N__35196;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35184;
    wire N__35181;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35169;
    wire N__35166;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35154;
    wire N__35151;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35139;
    wire N__35136;
    wire N__35135;
    wire N__35132;
    wire N__35129;
    wire N__35124;
    wire N__35121;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35109;
    wire N__35106;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35087;
    wire N__35086;
    wire N__35085;
    wire N__35084;
    wire N__35083;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35071;
    wire N__35064;
    wire N__35061;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35037;
    wire N__35036;
    wire N__35035;
    wire N__35032;
    wire N__35027;
    wire N__35022;
    wire N__35021;
    wire N__35018;
    wire N__35017;
    wire N__35014;
    wire N__35009;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34961;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34946;
    wire N__34943;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34916;
    wire N__34915;
    wire N__34914;
    wire N__34911;
    wire N__34910;
    wire N__34907;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34888;
    wire N__34887;
    wire N__34884;
    wire N__34879;
    wire N__34876;
    wire N__34869;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34856;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34839;
    wire N__34838;
    wire N__34837;
    wire N__34836;
    wire N__34833;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34815;
    wire N__34814;
    wire N__34813;
    wire N__34812;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34778;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34751;
    wire N__34746;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34727;
    wire N__34726;
    wire N__34723;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34439;
    wire N__34436;
    wire N__34431;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34421;
    wire N__34416;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34346;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34289;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34275;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34254;
    wire N__34251;
    wire N__34250;
    wire N__34247;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34224;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34212;
    wire N__34209;
    wire N__34208;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34176;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34142;
    wire N__34139;
    wire N__34138;
    wire N__34135;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34085;
    wire N__34082;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33959;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33944;
    wire N__33943;
    wire N__33942;
    wire N__33939;
    wire N__33932;
    wire N__33927;
    wire N__33924;
    wire N__33923;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33900;
    wire N__33897;
    wire N__33894;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33876;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33868;
    wire N__33861;
    wire N__33858;
    wire N__33857;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33845;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33833;
    wire N__33830;
    wire N__33829;
    wire N__33828;
    wire N__33825;
    wire N__33822;
    wire N__33817;
    wire N__33810;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33749;
    wire N__33748;
    wire N__33747;
    wire N__33744;
    wire N__33739;
    wire N__33736;
    wire N__33729;
    wire N__33726;
    wire N__33725;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33708;
    wire N__33707;
    wire N__33702;
    wire N__33699;
    wire N__33698;
    wire N__33697;
    wire N__33696;
    wire N__33695;
    wire N__33694;
    wire N__33693;
    wire N__33692;
    wire N__33691;
    wire N__33690;
    wire N__33689;
    wire N__33688;
    wire N__33687;
    wire N__33686;
    wire N__33685;
    wire N__33684;
    wire N__33683;
    wire N__33682;
    wire N__33681;
    wire N__33680;
    wire N__33679;
    wire N__33678;
    wire N__33677;
    wire N__33676;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33672;
    wire N__33671;
    wire N__33670;
    wire N__33669;
    wire N__33668;
    wire N__33659;
    wire N__33650;
    wire N__33643;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33619;
    wire N__33612;
    wire N__33603;
    wire N__33594;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33573;
    wire N__33562;
    wire N__33559;
    wire N__33552;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33497;
    wire N__33496;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33484;
    wire N__33481;
    wire N__33474;
    wire N__33473;
    wire N__33470;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33453;
    wire N__33452;
    wire N__33451;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33342;
    wire N__33341;
    wire N__33340;
    wire N__33339;
    wire N__33338;
    wire N__33337;
    wire N__33336;
    wire N__33335;
    wire N__33334;
    wire N__33333;
    wire N__33332;
    wire N__33331;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33282;
    wire N__33281;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33264;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33239;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33203;
    wire N__33202;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33159;
    wire N__33156;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33148;
    wire N__33143;
    wire N__33140;
    wire N__33137;
    wire N__33132;
    wire N__33129;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33119;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33107;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33037;
    wire N__33034;
    wire N__33027;
    wire N__33026;
    wire N__33023;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33008;
    wire N__33005;
    wire N__33000;
    wire N__32999;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32982;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32970;
    wire N__32967;
    wire N__32966;
    wire N__32963;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32947;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32915;
    wire N__32914;
    wire N__32911;
    wire N__32906;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32888;
    wire N__32887;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32858;
    wire N__32855;
    wire N__32854;
    wire N__32851;
    wire N__32848;
    wire N__32847;
    wire N__32844;
    wire N__32839;
    wire N__32836;
    wire N__32829;
    wire N__32828;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32801;
    wire N__32798;
    wire N__32797;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32772;
    wire N__32771;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32745;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32737;
    wire N__32734;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32691;
    wire N__32688;
    wire N__32685;
    wire N__32684;
    wire N__32683;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32646;
    wire N__32643;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32623;
    wire N__32616;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32605;
    wire N__32604;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32590;
    wire N__32583;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32559;
    wire N__32556;
    wire N__32555;
    wire N__32552;
    wire N__32551;
    wire N__32550;
    wire N__32545;
    wire N__32540;
    wire N__32535;
    wire N__32534;
    wire N__32533;
    wire N__32528;
    wire N__32527;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32515;
    wire N__32508;
    wire N__32507;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32490;
    wire N__32487;
    wire N__32486;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32471;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32453;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32387;
    wire N__32384;
    wire N__32381;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32006;
    wire N__32005;
    wire N__32002;
    wire N__31997;
    wire N__31992;
    wire N__31989;
    wire N__31988;
    wire N__31985;
    wire N__31984;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31958;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31946;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31934;
    wire N__31933;
    wire N__31930;
    wire N__31925;
    wire N__31920;
    wire N__31919;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31886;
    wire N__31883;
    wire N__31882;
    wire N__31877;
    wire N__31874;
    wire N__31871;
    wire N__31866;
    wire N__31863;
    wire N__31862;
    wire N__31861;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31845;
    wire N__31842;
    wire N__31841;
    wire N__31840;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31824;
    wire N__31821;
    wire N__31820;
    wire N__31817;
    wire N__31816;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31800;
    wire N__31797;
    wire N__31796;
    wire N__31793;
    wire N__31792;
    wire N__31787;
    wire N__31784;
    wire N__31781;
    wire N__31776;
    wire N__31773;
    wire N__31772;
    wire N__31771;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31755;
    wire N__31752;
    wire N__31751;
    wire N__31746;
    wire N__31745;
    wire N__31742;
    wire N__31739;
    wire N__31736;
    wire N__31731;
    wire N__31728;
    wire N__31727;
    wire N__31724;
    wire N__31719;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31704;
    wire N__31701;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31689;
    wire N__31686;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31674;
    wire N__31671;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31659;
    wire N__31656;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31644;
    wire N__31641;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31629;
    wire N__31626;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31614;
    wire N__31611;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31592;
    wire N__31591;
    wire N__31588;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31576;
    wire N__31571;
    wire N__31568;
    wire N__31563;
    wire N__31560;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31524;
    wire N__31521;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31509;
    wire N__31506;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31494;
    wire N__31491;
    wire N__31490;
    wire N__31487;
    wire N__31484;
    wire N__31479;
    wire N__31476;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31464;
    wire N__31461;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31449;
    wire N__31446;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31434;
    wire N__31431;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31419;
    wire N__31418;
    wire N__31415;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31397;
    wire N__31392;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31380;
    wire N__31377;
    wire N__31376;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31361;
    wire N__31356;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31338;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31307;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31265;
    wire N__31264;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31256;
    wire N__31255;
    wire N__31254;
    wire N__31251;
    wire N__31250;
    wire N__31249;
    wire N__31248;
    wire N__31245;
    wire N__31240;
    wire N__31239;
    wire N__31238;
    wire N__31237;
    wire N__31236;
    wire N__31235;
    wire N__31234;
    wire N__31233;
    wire N__31232;
    wire N__31231;
    wire N__31230;
    wire N__31229;
    wire N__31228;
    wire N__31227;
    wire N__31226;
    wire N__31225;
    wire N__31224;
    wire N__31223;
    wire N__31220;
    wire N__31219;
    wire N__31218;
    wire N__31217;
    wire N__31216;
    wire N__31215;
    wire N__31214;
    wire N__31213;
    wire N__31212;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31202;
    wire N__31201;
    wire N__31200;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31185;
    wire N__31178;
    wire N__31169;
    wire N__31166;
    wire N__31157;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31133;
    wire N__31124;
    wire N__31123;
    wire N__31122;
    wire N__31121;
    wire N__31120;
    wire N__31119;
    wire N__31118;
    wire N__31117;
    wire N__31114;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31092;
    wire N__31083;
    wire N__31080;
    wire N__31075;
    wire N__31068;
    wire N__31065;
    wire N__31058;
    wire N__31049;
    wire N__31038;
    wire N__31031;
    wire N__31026;
    wire N__31021;
    wire N__31014;
    wire N__31005;
    wire N__31004;
    wire N__31001;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30978;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30960;
    wire N__30953;
    wire N__30950;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30938;
    wire N__30935;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30920;
    wire N__30917;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30894;
    wire N__30893;
    wire N__30890;
    wire N__30889;
    wire N__30886;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30868;
    wire N__30863;
    wire N__30858;
    wire N__30857;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30836;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30824;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30777;
    wire N__30774;
    wire N__30773;
    wire N__30770;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30753;
    wire N__30752;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30744;
    wire N__30741;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30727;
    wire N__30724;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30669;
    wire N__30666;
    wire N__30663;
    wire N__30660;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30650;
    wire N__30647;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30632;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30611;
    wire N__30606;
    wire N__30605;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30566;
    wire N__30561;
    wire N__30560;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30299;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30284;
    wire N__30279;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30264;
    wire N__30261;
    wire N__30256;
    wire N__30253;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30228;
    wire N__30227;
    wire N__30224;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30213;
    wire N__30210;
    wire N__30205;
    wire N__30202;
    wire N__30197;
    wire N__30194;
    wire N__30189;
    wire N__30186;
    wire N__30185;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30162;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30154;
    wire N__30149;
    wire N__30146;
    wire N__30145;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30126;
    wire N__30125;
    wire N__30122;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30105;
    wire N__30104;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30087;
    wire N__30084;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30076;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29948;
    wire N__29943;
    wire N__29940;
    wire N__29939;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29927;
    wire N__29922;
    wire N__29921;
    wire N__29918;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29901;
    wire N__29898;
    wire N__29895;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29885;
    wire N__29882;
    wire N__29879;
    wire N__29874;
    wire N__29873;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29786;
    wire N__29785;
    wire N__29784;
    wire N__29783;
    wire N__29782;
    wire N__29779;
    wire N__29768;
    wire N__29765;
    wire N__29764;
    wire N__29763;
    wire N__29762;
    wire N__29759;
    wire N__29758;
    wire N__29755;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29737;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29658;
    wire N__29655;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29568;
    wire N__29565;
    wire N__29564;
    wire N__29561;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29531;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29472;
    wire N__29469;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29448;
    wire N__29445;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29432;
    wire N__29429;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29307;
    wire N__29304;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29243;
    wire N__29240;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29072;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29013;
    wire N__29010;
    wire N__29009;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28977;
    wire N__28974;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28966;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28917;
    wire N__28916;
    wire N__28911;
    wire N__28910;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28866;
    wire N__28865;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28842;
    wire N__28841;
    wire N__28840;
    wire N__28835;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28820;
    wire N__28815;
    wire N__28812;
    wire N__28811;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28799;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28776;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28758;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28668;
    wire N__28665;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28631;
    wire N__28628;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28611;
    wire N__28610;
    wire N__28609;
    wire N__28606;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28580;
    wire N__28575;
    wire N__28572;
    wire N__28571;
    wire N__28566;
    wire N__28563;
    wire N__28562;
    wire N__28559;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28542;
    wire N__28541;
    wire N__28540;
    wire N__28537;
    wire N__28536;
    wire N__28533;
    wire N__28528;
    wire N__28525;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28509;
    wire N__28508;
    wire N__28505;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28482;
    wire N__28481;
    wire N__28478;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28446;
    wire N__28445;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28423;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28402;
    wire N__28395;
    wire N__28394;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28364;
    wire N__28363;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28351;
    wire N__28344;
    wire N__28343;
    wire N__28340;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28323;
    wire N__28320;
    wire N__28319;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28280;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28265;
    wire N__28264;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28248;
    wire N__28245;
    wire N__28244;
    wire N__28243;
    wire N__28240;
    wire N__28235;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28220;
    wire N__28217;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28193;
    wire N__28190;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28160;
    wire N__28159;
    wire N__28156;
    wire N__28151;
    wire N__28146;
    wire N__28145;
    wire N__28142;
    wire N__28141;
    wire N__28138;
    wire N__28133;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28080;
    wire N__28077;
    wire N__28076;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28061;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28049;
    wire N__28048;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28032;
    wire N__28029;
    wire N__28028;
    wire N__28025;
    wire N__28024;
    wire N__28021;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28005;
    wire N__28002;
    wire N__28001;
    wire N__28000;
    wire N__27997;
    wire N__27992;
    wire N__27987;
    wire N__27984;
    wire N__27983;
    wire N__27982;
    wire N__27979;
    wire N__27974;
    wire N__27969;
    wire N__27966;
    wire N__27965;
    wire N__27964;
    wire N__27961;
    wire N__27956;
    wire N__27951;
    wire N__27948;
    wire N__27947;
    wire N__27946;
    wire N__27943;
    wire N__27938;
    wire N__27933;
    wire N__27930;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27915;
    wire N__27912;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27897;
    wire N__27894;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27879;
    wire N__27876;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27819;
    wire N__27816;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27762;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27747;
    wire N__27744;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27729;
    wire N__27726;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27711;
    wire N__27708;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27693;
    wire N__27690;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27680;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27654;
    wire N__27651;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27629;
    wire N__27626;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27609;
    wire N__27608;
    wire N__27605;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27588;
    wire N__27587;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27567;
    wire N__27564;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27543;
    wire N__27542;
    wire N__27539;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27522;
    wire N__27521;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27501;
    wire N__27500;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27480;
    wire N__27477;
    wire N__27476;
    wire N__27475;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27449;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27429;
    wire N__27426;
    wire N__27425;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27405;
    wire N__27404;
    wire N__27403;
    wire N__27402;
    wire N__27393;
    wire N__27392;
    wire N__27391;
    wire N__27390;
    wire N__27389;
    wire N__27388;
    wire N__27387;
    wire N__27384;
    wire N__27379;
    wire N__27370;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27173;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27158;
    wire N__27153;
    wire N__27150;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27135;
    wire N__27132;
    wire N__27131;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27116;
    wire N__27111;
    wire N__27108;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27093;
    wire N__27090;
    wire N__27089;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27074;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27062;
    wire N__27061;
    wire N__27060;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27015;
    wire N__27006;
    wire N__27005;
    wire N__27004;
    wire N__27003;
    wire N__27002;
    wire N__26991;
    wire N__26990;
    wire N__26989;
    wire N__26988;
    wire N__26985;
    wire N__26984;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26952;
    wire N__26949;
    wire N__26944;
    wire N__26941;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26918;
    wire N__26917;
    wire N__26916;
    wire N__26915;
    wire N__26914;
    wire N__26913;
    wire N__26912;
    wire N__26911;
    wire N__26908;
    wire N__26903;
    wire N__26900;
    wire N__26889;
    wire N__26884;
    wire N__26879;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26804;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26789;
    wire N__26784;
    wire N__26781;
    wire N__26780;
    wire N__26779;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26763;
    wire N__26760;
    wire N__26759;
    wire N__26758;
    wire N__26753;
    wire N__26750;
    wire N__26747;
    wire N__26742;
    wire N__26741;
    wire N__26740;
    wire N__26737;
    wire N__26732;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26698;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26682;
    wire N__26681;
    wire N__26678;
    wire N__26677;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26654;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26631;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26616;
    wire N__26613;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26605;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26589;
    wire N__26588;
    wire N__26587;
    wire N__26584;
    wire N__26579;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26545;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26522;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26507;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26492;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26462;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26447;
    wire N__26442;
    wire N__26439;
    wire N__26438;
    wire N__26433;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26418;
    wire N__26415;
    wire N__26414;
    wire N__26413;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26397;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26379;
    wire N__26376;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26360;
    wire N__26355;
    wire N__26352;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26344;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26328;
    wire N__26325;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26313;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26291;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26281;
    wire N__26276;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26264;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26249;
    wire N__26244;
    wire N__26241;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26230;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26214;
    wire N__26211;
    wire N__26210;
    wire N__26205;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26190;
    wire N__26187;
    wire N__26186;
    wire N__26185;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26169;
    wire N__26166;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26158;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26142;
    wire N__26141;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26126;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26109;
    wire N__26106;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26098;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26075;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26060;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26041;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__26018;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26003;
    wire N__25998;
    wire N__25995;
    wire N__25994;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25963;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25921;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25889;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25874;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25857;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25844;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25799;
    wire N__25794;
    wire N__25791;
    wire N__25790;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25764;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25695;
    wire N__25692;
    wire N__25691;
    wire N__25686;
    wire N__25683;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25617;
    wire N__25614;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25313;
    wire N__25312;
    wire N__25311;
    wire N__25308;
    wire N__25301;
    wire N__25296;
    wire N__25293;
    wire N__25292;
    wire N__25291;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25275;
    wire N__25274;
    wire N__25273;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25255;
    wire N__25248;
    wire N__25247;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25197;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25160;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25149;
    wire N__25146;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25122;
    wire N__25121;
    wire N__25120;
    wire N__25119;
    wire N__25118;
    wire N__25117;
    wire N__25116;
    wire N__25115;
    wire N__25114;
    wire N__25113;
    wire N__25112;
    wire N__25111;
    wire N__25110;
    wire N__25109;
    wire N__25108;
    wire N__25107;
    wire N__25106;
    wire N__25105;
    wire N__25104;
    wire N__25103;
    wire N__25102;
    wire N__25101;
    wire N__25100;
    wire N__25099;
    wire N__25098;
    wire N__25097;
    wire N__25096;
    wire N__25095;
    wire N__25094;
    wire N__25093;
    wire N__25084;
    wire N__25075;
    wire N__25066;
    wire N__25057;
    wire N__25048;
    wire N__25039;
    wire N__25034;
    wire N__25025;
    wire N__25012;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24932;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24917;
    wire N__24914;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24897;
    wire N__24896;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24873;
    wire N__24872;
    wire N__24867;
    wire N__24864;
    wire N__24863;
    wire N__24860;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24848;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24825;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24813;
    wire N__24810;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24770;
    wire N__24767;
    wire N__24766;
    wire N__24765;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24757;
    wire N__24756;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24738;
    wire N__24737;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24721;
    wire N__24718;
    wire N__24713;
    wire N__24706;
    wire N__24697;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24189;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24122;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24106;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24065;
    wire N__24062;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23966;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23943;
    wire N__23940;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23897;
    wire N__23894;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23754;
    wire N__23751;
    wire N__23750;
    wire N__23747;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23718;
    wire N__23715;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23597;
    wire N__23594;
    wire N__23593;
    wire N__23592;
    wire N__23591;
    wire N__23590;
    wire N__23589;
    wire N__23588;
    wire N__23587;
    wire N__23586;
    wire N__23585;
    wire N__23584;
    wire N__23583;
    wire N__23582;
    wire N__23581;
    wire N__23580;
    wire N__23579;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23556;
    wire N__23553;
    wire N__23552;
    wire N__23549;
    wire N__23534;
    wire N__23531;
    wire N__23530;
    wire N__23529;
    wire N__23528;
    wire N__23527;
    wire N__23526;
    wire N__23525;
    wire N__23524;
    wire N__23523;
    wire N__23522;
    wire N__23521;
    wire N__23520;
    wire N__23519;
    wire N__23510;
    wire N__23507;
    wire N__23506;
    wire N__23501;
    wire N__23498;
    wire N__23491;
    wire N__23488;
    wire N__23477;
    wire N__23474;
    wire N__23463;
    wire N__23458;
    wire N__23455;
    wire N__23450;
    wire N__23445;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23427;
    wire N__23426;
    wire N__23425;
    wire N__23424;
    wire N__23423;
    wire N__23422;
    wire N__23421;
    wire N__23420;
    wire N__23419;
    wire N__23418;
    wire N__23417;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23391;
    wire N__23390;
    wire N__23389;
    wire N__23388;
    wire N__23387;
    wire N__23382;
    wire N__23381;
    wire N__23380;
    wire N__23379;
    wire N__23378;
    wire N__23375;
    wire N__23374;
    wire N__23373;
    wire N__23372;
    wire N__23371;
    wire N__23370;
    wire N__23369;
    wire N__23366;
    wire N__23359;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23341;
    wire N__23340;
    wire N__23339;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23305;
    wire N__23300;
    wire N__23289;
    wire N__23284;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23246;
    wire N__23245;
    wire N__23244;
    wire N__23243;
    wire N__23242;
    wire N__23241;
    wire N__23240;
    wire N__23239;
    wire N__23238;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23223;
    wire N__23222;
    wire N__23221;
    wire N__23218;
    wire N__23217;
    wire N__23214;
    wire N__23213;
    wire N__23212;
    wire N__23209;
    wire N__23208;
    wire N__23207;
    wire N__23206;
    wire N__23205;
    wire N__23204;
    wire N__23203;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23197;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23182;
    wire N__23179;
    wire N__23172;
    wire N__23167;
    wire N__23164;
    wire N__23159;
    wire N__23152;
    wire N__23151;
    wire N__23150;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23126;
    wire N__23123;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23096;
    wire N__23093;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23067;
    wire N__23062;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23012;
    wire N__23009;
    wire N__23008;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22987;
    wire N__22984;
    wire N__22977;
    wire N__22974;
    wire N__22973;
    wire N__22970;
    wire N__22969;
    wire N__22966;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22946;
    wire N__22943;
    wire N__22938;
    wire N__22935;
    wire N__22934;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22917;
    wire N__22914;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22883;
    wire N__22882;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22853;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22811;
    wire N__22810;
    wire N__22805;
    wire N__22802;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22784;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22769;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22757;
    wire N__22756;
    wire N__22751;
    wire N__22748;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22718;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22697;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22670;
    wire N__22669;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22595;
    wire N__22594;
    wire N__22591;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22563;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22488;
    wire N__22485;
    wire N__22484;
    wire N__22481;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22463;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22448;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22415;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22316;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22275;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22240;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22219;
    wire N__22216;
    wire N__22209;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22197;
    wire N__22194;
    wire N__22191;
    wire N__22190;
    wire N__22187;
    wire N__22186;
    wire N__22183;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22165;
    wire N__22162;
    wire N__22155;
    wire N__22154;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22136;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22104;
    wire N__22101;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22076;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22068;
    wire N__22065;
    wire N__22060;
    wire N__22057;
    wire N__22050;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22019;
    wire N__22018;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22000;
    wire N__21997;
    wire N__21990;
    wire N__21989;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21974;
    wire N__21971;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21936;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21908;
    wire N__21907;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21895;
    wire N__21888;
    wire N__21887;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21872;
    wire N__21869;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21858;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21840;
    wire N__21839;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21779;
    wire N__21778;
    wire N__21775;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21757;
    wire N__21750;
    wire N__21749;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21719;
    wire N__21718;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21700;
    wire N__21693;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21674;
    wire N__21671;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21646;
    wire N__21639;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21620;
    wire N__21619;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21588;
    wire N__21585;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21559;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21541;
    wire N__21538;
    wire N__21531;
    wire N__21530;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21509;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21495;
    wire N__21492;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21474;
    wire N__21471;
    wire N__21470;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21453;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21435;
    wire N__21432;
    wire N__21431;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21401;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21380;
    wire N__21377;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21366;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21350;
    wire N__21347;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21329;
    wire N__21326;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21311;
    wire N__21308;
    wire N__21307;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21289;
    wire N__21286;
    wire N__21279;
    wire N__21278;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21257;
    wire N__21254;
    wire N__21253;
    wire N__21250;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21210;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21198;
    wire N__21195;
    wire N__21194;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21141;
    wire N__21138;
    wire N__21137;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21017;
    wire N__21016;
    wire N__21013;
    wire N__21012;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20975;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20930;
    wire N__20929;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20895;
    wire N__20894;
    wire N__20891;
    wire N__20890;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20875;
    wire N__20872;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20633;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20613;
    wire N__20612;
    wire N__20609;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20594;
    wire N__20589;
    wire N__20588;
    wire N__20585;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20565;
    wire N__20562;
    wire N__20561;
    wire N__20560;
    wire N__20557;
    wire N__20552;
    wire N__20549;
    wire N__20544;
    wire N__20543;
    wire N__20542;
    wire N__20539;
    wire N__20534;
    wire N__20531;
    wire N__20526;
    wire N__20525;
    wire N__20524;
    wire N__20521;
    wire N__20516;
    wire N__20513;
    wire N__20508;
    wire N__20505;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20483;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20375;
    wire N__20374;
    wire N__20373;
    wire N__20372;
    wire N__20371;
    wire N__20370;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20333;
    wire N__20332;
    wire N__20325;
    wire N__20322;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20310;
    wire N__20309;
    wire N__20304;
    wire N__20301;
    wire N__20300;
    wire N__20299;
    wire N__20296;
    wire N__20295;
    wire N__20294;
    wire N__20289;
    wire N__20282;
    wire N__20281;
    wire N__20280;
    wire N__20275;
    wire N__20274;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20232;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20211;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19241;
    wire N__19240;
    wire N__19239;
    wire N__19238;
    wire N__19237;
    wire N__19236;
    wire N__19235;
    wire N__19234;
    wire N__19233;
    wire N__19232;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19185;
    wire N__19176;
    wire N__19171;
    wire N__19166;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19077;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_1_9_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_1_10_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire bfn_1_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire bfn_1_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire bfn_1_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire bfn_1_15_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire un7_start_stop;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44 ;
    wire \current_shift_inst.PI_CTRL.N_77 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.N_43_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_98_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_158 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.N_96_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_160 ;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire pwm_duty_input_0;
    wire \pwm_generator_inst.un2_duty_input_0_o3_1Z0Z_0 ;
    wire \pwm_generator_inst.N_7_cascade_ ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_6;
    wire pwm_duty_input_7;
    wire pwm_duty_input_8;
    wire pwm_duty_input_3;
    wire pwm_duty_input_4;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_2_24_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_2_25_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire bfn_2_26_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire N_88_i_i;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire bfn_3_17_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire bfn_3_18_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire bfn_3_19_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire bfn_3_20_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire bfn_3_24_0_;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire bfn_3_25_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.N_46 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire bfn_4_22_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire bfn_4_23_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire bfn_4_24_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_30 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire bfn_5_23_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire bfn_5_24_0_;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire bfn_5_25_0_;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire bfn_7_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_7_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_7_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_7_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_166_i ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ;
    wire bfn_7_26_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_7_27_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_8_1_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_8_2_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire bfn_8_3_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire elapsed_time_ns_1_RNI0BPBB_0_22_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire elapsed_time_ns_1_RNI3EPBB_0_25_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_8_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire bfn_8_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_8_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_8_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_165_i ;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_8_24_0_;
    wire \pwm_generator_inst.threshold_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.threshold_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.threshold_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.threshold_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_8_25_0_;
    wire \pwm_generator_inst.threshold_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_9_3_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_9_4_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_9_5_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_9_6_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_9_13_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire bfn_9_14_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire bfn_9_15_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire bfn_9_16_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_27 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_28 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_30 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_10_8_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_10_9_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire bfn_10_10_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire elapsed_time_ns_1_RNI1BOBB_0_14_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire bfn_11_8_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_11_10_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_11_11_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \current_shift_inst.N_1263_i ;
    wire \current_shift_inst.control_input_1 ;
    wire bfn_11_13_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_11_14_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.control_input_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire \current_shift_inst.control_input_cry_14 ;
    wire \current_shift_inst.control_input_cry_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire bfn_11_15_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.control_input_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.control_input_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.control_input_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.control_input_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.control_input_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.control_input_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.control_input_cry_22 ;
    wire \current_shift_inst.control_input_cry_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.control_input_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ;
    wire \current_shift_inst.control_input_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ;
    wire \current_shift_inst.control_input_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ;
    wire \current_shift_inst.control_input_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ;
    wire \current_shift_inst.control_input_cry_28 ;
    wire \current_shift_inst.control_input_cry_29 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.control_input_axb_26 ;
    wire \current_shift_inst.control_input_axb_29 ;
    wire \current_shift_inst.control_input_axb_17 ;
    wire s4_phy_c;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire il_max_comp2_c;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.N_54_0 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.control_input_axb_13 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.control_input_axb_15 ;
    wire \current_shift_inst.control_input_axb_14 ;
    wire \current_shift_inst.control_input_axb_16 ;
    wire \current_shift_inst.control_input_axb_18 ;
    wire \current_shift_inst.control_input_axb_19 ;
    wire \current_shift_inst.control_input_axb_20 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.control_input_axb_23 ;
    wire \current_shift_inst.control_input_axb_24 ;
    wire \current_shift_inst.control_input_axb_25 ;
    wire \current_shift_inst.control_input_axb_27 ;
    wire delay_hc_input_c_g;
    wire s3_phy_c;
    wire GB_BUFFER_red_c_g_THRU_CO;
    wire \phase_controller_inst1.state_ns_0_0_1 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.start_flagZ0 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.N_54_0 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire il_max_comp1_c;
    wire \phase_controller_inst2.state_ns_0_0_1 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.N_61 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_13_8_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_13_9_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire bfn_13_10_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire elapsed_time_ns_1_RNII43T9_0_6_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire elapsed_time_ns_1_RNI69DN9_0_28_cascade_;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire bfn_13_16_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire bfn_13_17_0_;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire bfn_13_18_0_;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire bfn_13_19_0_;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire s2_phy_c;
    wire state_3;
    wire s1_phy_c;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_161_i ;
    wire il_min_comp1_c;
    wire \phase_controller_inst1.N_61 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire start_stop_c;
    wire \phase_controller_inst2.stateZ0Z_4 ;
    wire \phase_controller_inst2.start_flagZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_14_7_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_14_8_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_14_9_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_14_10_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire bfn_14_13_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire bfn_14_14_0_;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.control_input_axb_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire \current_shift_inst.control_input_axb_21 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_0_s0_4 ;
    wire \current_shift_inst.un38_control_input_0_s1_4 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.un38_control_input_0_s0_3 ;
    wire \current_shift_inst.un38_control_input_0_s1_3 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire bfn_15_21_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_15_22_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_15_23_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_15_24_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_16_7_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_16_8_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire bfn_16_9_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire bfn_16_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire bfn_16_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire bfn_16_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_16_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_16_19_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_16_20_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_16_21_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_16_22_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_17_7_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_17_8_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_17_9_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_17_10_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ;
    wire bfn_17_15_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_17_16_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire bfn_17_17_0_;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire bfn_17_23_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_17_24_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_17_25_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_17_26_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_162_i ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire bfn_18_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_18_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_18_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_18_14_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.N_161_i_g ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.N_164_i ;
    wire \delay_measurement_inst.delay_hc_timer.N_163_i ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire clk_100mhz_0;
    wire red_c_g;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire N_19_1;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__27351),
            .RESETB(N__33516),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38709),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38706),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__29838,N__29861,N__29499,N__29532,N__29565,N__29598,N__29624,N__29654,N__29685,N__29711,N__29270,N__29304,N__29334,N__29358,N__29391,N__29415}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__38708,dangling_wire_45,N__38707}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38862),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38855),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__48866,N__48859,N__48864,N__48858,N__48865,N__48857,N__48867,N__48854,N__48860,N__48853,N__48861,N__48855,N__48862,N__48856,N__48863}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__38861,N__38858,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__38856,N__38860,N__38857,N__38859}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38677),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38670),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__48835,N__48838,N__48836,N__48839,N__48837,N__20634,N__20565,N__20588,N__20613,N__20504,N__20526,N__20544,N__20232,N__20247,N__20211}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__38676,N__38673,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__38671,N__38675,N__38672,N__38674}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38758),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38755),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__29445,N__29469,N__29010,N__29043,N__29076,N__29106,N__29139,N__29169,N__29193,N__29214,N__29243,N__28665,N__28695,N__28733,N__30807}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__38757,dangling_wire_215,N__38756}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__50509),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__50511),
            .DIN(N__50510),
            .DOUT(N__50509),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__50511),
            .PADOUT(N__50510),
            .PADIN(N__50509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__50500),
            .DIN(N__50499),
            .DOUT(N__50498),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__50500),
            .PADOUT(N__50499),
            .PADIN(N__50498),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__50491),
            .DIN(N__50490),
            .DOUT(N__50489),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__50491),
            .PADOUT(N__50490),
            .PADIN(N__50489),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__50482),
            .DIN(N__50481),
            .DOUT(N__50480),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__50482),
            .PADOUT(N__50481),
            .PADIN(N__50480),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27201),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__50473),
            .DIN(N__50472),
            .DOUT(N__50471),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__50473),
            .PADOUT(N__50472),
            .PADIN(N__50471),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__50464),
            .DIN(N__50463),
            .DOUT(N__50462),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__50464),
            .PADOUT(N__50463),
            .PADIN(N__50462),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34926),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__50455),
            .DIN(N__50454),
            .DOUT(N__50453),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__50455),
            .PADOUT(N__50454),
            .PADIN(N__50453),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__50446),
            .DIN(N__50445),
            .DOUT(N__50444),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__50446),
            .PADOUT(N__50445),
            .PADIN(N__50444),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34869),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__50437),
            .DIN(N__50436),
            .DOUT(N__50435),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__50437),
            .PADOUT(N__50436),
            .PADIN(N__50435),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32355),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__50428),
            .DIN(N__50427),
            .DOUT(N__50426),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__50428),
            .PADOUT(N__50427),
            .PADIN(N__50426),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__50419),
            .DIN(N__50418),
            .DOUT(N__50417),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__50419),
            .PADOUT(N__50418),
            .PADIN(N__50417),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33534),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__50410),
            .DIN(N__50409),
            .DOUT(N__50408),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__50410),
            .PADOUT(N__50409),
            .PADIN(N__50408),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__50401),
            .DIN(N__50400),
            .DOUT(N__50399),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__50401),
            .PADOUT(N__50400),
            .PADIN(N__50399),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__12029 (
            .O(N__50382),
            .I(N__50379));
    LocalMux I__12028 (
            .O(N__50379),
            .I(N__50376));
    Span4Mux_v I__12027 (
            .O(N__50376),
            .I(N__50372));
    InMux I__12026 (
            .O(N__50375),
            .I(N__50368));
    Span4Mux_h I__12025 (
            .O(N__50372),
            .I(N__50365));
    InMux I__12024 (
            .O(N__50371),
            .I(N__50362));
    LocalMux I__12023 (
            .O(N__50368),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__12022 (
            .O(N__50365),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    LocalMux I__12021 (
            .O(N__50362),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    CascadeMux I__12020 (
            .O(N__50355),
            .I(N__50352));
    InMux I__12019 (
            .O(N__50352),
            .I(N__50348));
    InMux I__12018 (
            .O(N__50351),
            .I(N__50345));
    LocalMux I__12017 (
            .O(N__50348),
            .I(N__50341));
    LocalMux I__12016 (
            .O(N__50345),
            .I(N__50338));
    InMux I__12015 (
            .O(N__50344),
            .I(N__50335));
    Span4Mux_v I__12014 (
            .O(N__50341),
            .I(N__50332));
    Odrv4 I__12013 (
            .O(N__50338),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__12012 (
            .O(N__50335),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__12011 (
            .O(N__50332),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__12010 (
            .O(N__50325),
            .I(N__50320));
    InMux I__12009 (
            .O(N__50324),
            .I(N__50316));
    InMux I__12008 (
            .O(N__50323),
            .I(N__50313));
    LocalMux I__12007 (
            .O(N__50320),
            .I(N__50310));
    InMux I__12006 (
            .O(N__50319),
            .I(N__50307));
    LocalMux I__12005 (
            .O(N__50316),
            .I(N__50304));
    LocalMux I__12004 (
            .O(N__50313),
            .I(N__50301));
    Span4Mux_v I__12003 (
            .O(N__50310),
            .I(N__50296));
    LocalMux I__12002 (
            .O(N__50307),
            .I(N__50296));
    Span4Mux_h I__12001 (
            .O(N__50304),
            .I(N__50293));
    Span4Mux_v I__12000 (
            .O(N__50301),
            .I(N__50288));
    Span4Mux_h I__11999 (
            .O(N__50296),
            .I(N__50288));
    Odrv4 I__11998 (
            .O(N__50293),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__11997 (
            .O(N__50288),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    CEMux I__11996 (
            .O(N__50283),
            .I(N__50280));
    LocalMux I__11995 (
            .O(N__50280),
            .I(N__50274));
    CEMux I__11994 (
            .O(N__50279),
            .I(N__50271));
    CEMux I__11993 (
            .O(N__50278),
            .I(N__50268));
    CEMux I__11992 (
            .O(N__50277),
            .I(N__50265));
    Span4Mux_v I__11991 (
            .O(N__50274),
            .I(N__50260));
    LocalMux I__11990 (
            .O(N__50271),
            .I(N__50260));
    LocalMux I__11989 (
            .O(N__50268),
            .I(N__50257));
    LocalMux I__11988 (
            .O(N__50265),
            .I(N__50254));
    Span4Mux_v I__11987 (
            .O(N__50260),
            .I(N__50251));
    Span4Mux_h I__11986 (
            .O(N__50257),
            .I(N__50248));
    Span4Mux_h I__11985 (
            .O(N__50254),
            .I(N__50245));
    Odrv4 I__11984 (
            .O(N__50251),
            .I(\delay_measurement_inst.delay_hc_timer.N_164_i ));
    Odrv4 I__11983 (
            .O(N__50248),
            .I(\delay_measurement_inst.delay_hc_timer.N_164_i ));
    Odrv4 I__11982 (
            .O(N__50245),
            .I(\delay_measurement_inst.delay_hc_timer.N_164_i ));
    CEMux I__11981 (
            .O(N__50238),
            .I(N__50235));
    LocalMux I__11980 (
            .O(N__50235),
            .I(N__50230));
    CEMux I__11979 (
            .O(N__50234),
            .I(N__50227));
    CEMux I__11978 (
            .O(N__50233),
            .I(N__50223));
    Span4Mux_v I__11977 (
            .O(N__50230),
            .I(N__50218));
    LocalMux I__11976 (
            .O(N__50227),
            .I(N__50218));
    CEMux I__11975 (
            .O(N__50226),
            .I(N__50215));
    LocalMux I__11974 (
            .O(N__50223),
            .I(N__50211));
    Span4Mux_h I__11973 (
            .O(N__50218),
            .I(N__50208));
    LocalMux I__11972 (
            .O(N__50215),
            .I(N__50205));
    CEMux I__11971 (
            .O(N__50214),
            .I(N__50202));
    Span4Mux_h I__11970 (
            .O(N__50211),
            .I(N__50199));
    Span4Mux_h I__11969 (
            .O(N__50208),
            .I(N__50196));
    Span4Mux_h I__11968 (
            .O(N__50205),
            .I(N__50191));
    LocalMux I__11967 (
            .O(N__50202),
            .I(N__50191));
    Odrv4 I__11966 (
            .O(N__50199),
            .I(\delay_measurement_inst.delay_hc_timer.N_163_i ));
    Odrv4 I__11965 (
            .O(N__50196),
            .I(\delay_measurement_inst.delay_hc_timer.N_163_i ));
    Odrv4 I__11964 (
            .O(N__50191),
            .I(\delay_measurement_inst.delay_hc_timer.N_163_i ));
    InMux I__11963 (
            .O(N__50184),
            .I(N__50150));
    InMux I__11962 (
            .O(N__50183),
            .I(N__50150));
    InMux I__11961 (
            .O(N__50182),
            .I(N__50150));
    InMux I__11960 (
            .O(N__50181),
            .I(N__50150));
    InMux I__11959 (
            .O(N__50180),
            .I(N__50137));
    InMux I__11958 (
            .O(N__50179),
            .I(N__50137));
    InMux I__11957 (
            .O(N__50178),
            .I(N__50137));
    InMux I__11956 (
            .O(N__50177),
            .I(N__50137));
    InMux I__11955 (
            .O(N__50176),
            .I(N__50128));
    InMux I__11954 (
            .O(N__50175),
            .I(N__50128));
    InMux I__11953 (
            .O(N__50174),
            .I(N__50128));
    InMux I__11952 (
            .O(N__50173),
            .I(N__50128));
    InMux I__11951 (
            .O(N__50172),
            .I(N__50123));
    InMux I__11950 (
            .O(N__50171),
            .I(N__50123));
    InMux I__11949 (
            .O(N__50170),
            .I(N__50114));
    InMux I__11948 (
            .O(N__50169),
            .I(N__50114));
    InMux I__11947 (
            .O(N__50168),
            .I(N__50114));
    InMux I__11946 (
            .O(N__50167),
            .I(N__50114));
    InMux I__11945 (
            .O(N__50166),
            .I(N__50105));
    InMux I__11944 (
            .O(N__50165),
            .I(N__50105));
    InMux I__11943 (
            .O(N__50164),
            .I(N__50105));
    InMux I__11942 (
            .O(N__50163),
            .I(N__50105));
    InMux I__11941 (
            .O(N__50162),
            .I(N__50096));
    InMux I__11940 (
            .O(N__50161),
            .I(N__50096));
    InMux I__11939 (
            .O(N__50160),
            .I(N__50096));
    InMux I__11938 (
            .O(N__50159),
            .I(N__50096));
    LocalMux I__11937 (
            .O(N__50150),
            .I(N__50093));
    InMux I__11936 (
            .O(N__50149),
            .I(N__50084));
    InMux I__11935 (
            .O(N__50148),
            .I(N__50084));
    InMux I__11934 (
            .O(N__50147),
            .I(N__50084));
    InMux I__11933 (
            .O(N__50146),
            .I(N__50084));
    LocalMux I__11932 (
            .O(N__50137),
            .I(N__50079));
    LocalMux I__11931 (
            .O(N__50128),
            .I(N__50079));
    LocalMux I__11930 (
            .O(N__50123),
            .I(N__50076));
    LocalMux I__11929 (
            .O(N__50114),
            .I(N__50073));
    LocalMux I__11928 (
            .O(N__50105),
            .I(N__50068));
    LocalMux I__11927 (
            .O(N__50096),
            .I(N__50068));
    Span4Mux_v I__11926 (
            .O(N__50093),
            .I(N__50063));
    LocalMux I__11925 (
            .O(N__50084),
            .I(N__50063));
    Span4Mux_h I__11924 (
            .O(N__50079),
            .I(N__50060));
    Span4Mux_h I__11923 (
            .O(N__50076),
            .I(N__50055));
    Span4Mux_h I__11922 (
            .O(N__50073),
            .I(N__50055));
    Span4Mux_h I__11921 (
            .O(N__50068),
            .I(N__50052));
    Odrv4 I__11920 (
            .O(N__50063),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__11919 (
            .O(N__50060),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__11918 (
            .O(N__50055),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__11917 (
            .O(N__50052),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__11916 (
            .O(N__50043),
            .I(N__50039));
    CascadeMux I__11915 (
            .O(N__50042),
            .I(N__50036));
    LocalMux I__11914 (
            .O(N__50039),
            .I(N__50032));
    InMux I__11913 (
            .O(N__50036),
            .I(N__50027));
    InMux I__11912 (
            .O(N__50035),
            .I(N__50027));
    Span4Mux_v I__11911 (
            .O(N__50032),
            .I(N__50022));
    LocalMux I__11910 (
            .O(N__50027),
            .I(N__50022));
    Span4Mux_h I__11909 (
            .O(N__50022),
            .I(N__50019));
    Span4Mux_h I__11908 (
            .O(N__50019),
            .I(N__50016));
    Span4Mux_v I__11907 (
            .O(N__50016),
            .I(N__50013));
    Odrv4 I__11906 (
            .O(N__50013),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__11905 (
            .O(N__50010),
            .I(N__50007));
    LocalMux I__11904 (
            .O(N__50007),
            .I(N__50003));
    InMux I__11903 (
            .O(N__50006),
            .I(N__50000));
    Span4Mux_v I__11902 (
            .O(N__50003),
            .I(N__49995));
    LocalMux I__11901 (
            .O(N__50000),
            .I(N__49995));
    Span4Mux_h I__11900 (
            .O(N__49995),
            .I(N__49992));
    Span4Mux_h I__11899 (
            .O(N__49992),
            .I(N__49987));
    InMux I__11898 (
            .O(N__49991),
            .I(N__49982));
    InMux I__11897 (
            .O(N__49990),
            .I(N__49982));
    Span4Mux_v I__11896 (
            .O(N__49987),
            .I(N__49979));
    LocalMux I__11895 (
            .O(N__49982),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__11894 (
            .O(N__49979),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__11893 (
            .O(N__49974),
            .I(N__49968));
    InMux I__11892 (
            .O(N__49973),
            .I(N__49961));
    InMux I__11891 (
            .O(N__49972),
            .I(N__49961));
    InMux I__11890 (
            .O(N__49971),
            .I(N__49961));
    LocalMux I__11889 (
            .O(N__49968),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__11888 (
            .O(N__49961),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    ClkMux I__11887 (
            .O(N__49956),
            .I(N__49482));
    ClkMux I__11886 (
            .O(N__49955),
            .I(N__49482));
    ClkMux I__11885 (
            .O(N__49954),
            .I(N__49482));
    ClkMux I__11884 (
            .O(N__49953),
            .I(N__49482));
    ClkMux I__11883 (
            .O(N__49952),
            .I(N__49482));
    ClkMux I__11882 (
            .O(N__49951),
            .I(N__49482));
    ClkMux I__11881 (
            .O(N__49950),
            .I(N__49482));
    ClkMux I__11880 (
            .O(N__49949),
            .I(N__49482));
    ClkMux I__11879 (
            .O(N__49948),
            .I(N__49482));
    ClkMux I__11878 (
            .O(N__49947),
            .I(N__49482));
    ClkMux I__11877 (
            .O(N__49946),
            .I(N__49482));
    ClkMux I__11876 (
            .O(N__49945),
            .I(N__49482));
    ClkMux I__11875 (
            .O(N__49944),
            .I(N__49482));
    ClkMux I__11874 (
            .O(N__49943),
            .I(N__49482));
    ClkMux I__11873 (
            .O(N__49942),
            .I(N__49482));
    ClkMux I__11872 (
            .O(N__49941),
            .I(N__49482));
    ClkMux I__11871 (
            .O(N__49940),
            .I(N__49482));
    ClkMux I__11870 (
            .O(N__49939),
            .I(N__49482));
    ClkMux I__11869 (
            .O(N__49938),
            .I(N__49482));
    ClkMux I__11868 (
            .O(N__49937),
            .I(N__49482));
    ClkMux I__11867 (
            .O(N__49936),
            .I(N__49482));
    ClkMux I__11866 (
            .O(N__49935),
            .I(N__49482));
    ClkMux I__11865 (
            .O(N__49934),
            .I(N__49482));
    ClkMux I__11864 (
            .O(N__49933),
            .I(N__49482));
    ClkMux I__11863 (
            .O(N__49932),
            .I(N__49482));
    ClkMux I__11862 (
            .O(N__49931),
            .I(N__49482));
    ClkMux I__11861 (
            .O(N__49930),
            .I(N__49482));
    ClkMux I__11860 (
            .O(N__49929),
            .I(N__49482));
    ClkMux I__11859 (
            .O(N__49928),
            .I(N__49482));
    ClkMux I__11858 (
            .O(N__49927),
            .I(N__49482));
    ClkMux I__11857 (
            .O(N__49926),
            .I(N__49482));
    ClkMux I__11856 (
            .O(N__49925),
            .I(N__49482));
    ClkMux I__11855 (
            .O(N__49924),
            .I(N__49482));
    ClkMux I__11854 (
            .O(N__49923),
            .I(N__49482));
    ClkMux I__11853 (
            .O(N__49922),
            .I(N__49482));
    ClkMux I__11852 (
            .O(N__49921),
            .I(N__49482));
    ClkMux I__11851 (
            .O(N__49920),
            .I(N__49482));
    ClkMux I__11850 (
            .O(N__49919),
            .I(N__49482));
    ClkMux I__11849 (
            .O(N__49918),
            .I(N__49482));
    ClkMux I__11848 (
            .O(N__49917),
            .I(N__49482));
    ClkMux I__11847 (
            .O(N__49916),
            .I(N__49482));
    ClkMux I__11846 (
            .O(N__49915),
            .I(N__49482));
    ClkMux I__11845 (
            .O(N__49914),
            .I(N__49482));
    ClkMux I__11844 (
            .O(N__49913),
            .I(N__49482));
    ClkMux I__11843 (
            .O(N__49912),
            .I(N__49482));
    ClkMux I__11842 (
            .O(N__49911),
            .I(N__49482));
    ClkMux I__11841 (
            .O(N__49910),
            .I(N__49482));
    ClkMux I__11840 (
            .O(N__49909),
            .I(N__49482));
    ClkMux I__11839 (
            .O(N__49908),
            .I(N__49482));
    ClkMux I__11838 (
            .O(N__49907),
            .I(N__49482));
    ClkMux I__11837 (
            .O(N__49906),
            .I(N__49482));
    ClkMux I__11836 (
            .O(N__49905),
            .I(N__49482));
    ClkMux I__11835 (
            .O(N__49904),
            .I(N__49482));
    ClkMux I__11834 (
            .O(N__49903),
            .I(N__49482));
    ClkMux I__11833 (
            .O(N__49902),
            .I(N__49482));
    ClkMux I__11832 (
            .O(N__49901),
            .I(N__49482));
    ClkMux I__11831 (
            .O(N__49900),
            .I(N__49482));
    ClkMux I__11830 (
            .O(N__49899),
            .I(N__49482));
    ClkMux I__11829 (
            .O(N__49898),
            .I(N__49482));
    ClkMux I__11828 (
            .O(N__49897),
            .I(N__49482));
    ClkMux I__11827 (
            .O(N__49896),
            .I(N__49482));
    ClkMux I__11826 (
            .O(N__49895),
            .I(N__49482));
    ClkMux I__11825 (
            .O(N__49894),
            .I(N__49482));
    ClkMux I__11824 (
            .O(N__49893),
            .I(N__49482));
    ClkMux I__11823 (
            .O(N__49892),
            .I(N__49482));
    ClkMux I__11822 (
            .O(N__49891),
            .I(N__49482));
    ClkMux I__11821 (
            .O(N__49890),
            .I(N__49482));
    ClkMux I__11820 (
            .O(N__49889),
            .I(N__49482));
    ClkMux I__11819 (
            .O(N__49888),
            .I(N__49482));
    ClkMux I__11818 (
            .O(N__49887),
            .I(N__49482));
    ClkMux I__11817 (
            .O(N__49886),
            .I(N__49482));
    ClkMux I__11816 (
            .O(N__49885),
            .I(N__49482));
    ClkMux I__11815 (
            .O(N__49884),
            .I(N__49482));
    ClkMux I__11814 (
            .O(N__49883),
            .I(N__49482));
    ClkMux I__11813 (
            .O(N__49882),
            .I(N__49482));
    ClkMux I__11812 (
            .O(N__49881),
            .I(N__49482));
    ClkMux I__11811 (
            .O(N__49880),
            .I(N__49482));
    ClkMux I__11810 (
            .O(N__49879),
            .I(N__49482));
    ClkMux I__11809 (
            .O(N__49878),
            .I(N__49482));
    ClkMux I__11808 (
            .O(N__49877),
            .I(N__49482));
    ClkMux I__11807 (
            .O(N__49876),
            .I(N__49482));
    ClkMux I__11806 (
            .O(N__49875),
            .I(N__49482));
    ClkMux I__11805 (
            .O(N__49874),
            .I(N__49482));
    ClkMux I__11804 (
            .O(N__49873),
            .I(N__49482));
    ClkMux I__11803 (
            .O(N__49872),
            .I(N__49482));
    ClkMux I__11802 (
            .O(N__49871),
            .I(N__49482));
    ClkMux I__11801 (
            .O(N__49870),
            .I(N__49482));
    ClkMux I__11800 (
            .O(N__49869),
            .I(N__49482));
    ClkMux I__11799 (
            .O(N__49868),
            .I(N__49482));
    ClkMux I__11798 (
            .O(N__49867),
            .I(N__49482));
    ClkMux I__11797 (
            .O(N__49866),
            .I(N__49482));
    ClkMux I__11796 (
            .O(N__49865),
            .I(N__49482));
    ClkMux I__11795 (
            .O(N__49864),
            .I(N__49482));
    ClkMux I__11794 (
            .O(N__49863),
            .I(N__49482));
    ClkMux I__11793 (
            .O(N__49862),
            .I(N__49482));
    ClkMux I__11792 (
            .O(N__49861),
            .I(N__49482));
    ClkMux I__11791 (
            .O(N__49860),
            .I(N__49482));
    ClkMux I__11790 (
            .O(N__49859),
            .I(N__49482));
    ClkMux I__11789 (
            .O(N__49858),
            .I(N__49482));
    ClkMux I__11788 (
            .O(N__49857),
            .I(N__49482));
    ClkMux I__11787 (
            .O(N__49856),
            .I(N__49482));
    ClkMux I__11786 (
            .O(N__49855),
            .I(N__49482));
    ClkMux I__11785 (
            .O(N__49854),
            .I(N__49482));
    ClkMux I__11784 (
            .O(N__49853),
            .I(N__49482));
    ClkMux I__11783 (
            .O(N__49852),
            .I(N__49482));
    ClkMux I__11782 (
            .O(N__49851),
            .I(N__49482));
    ClkMux I__11781 (
            .O(N__49850),
            .I(N__49482));
    ClkMux I__11780 (
            .O(N__49849),
            .I(N__49482));
    ClkMux I__11779 (
            .O(N__49848),
            .I(N__49482));
    ClkMux I__11778 (
            .O(N__49847),
            .I(N__49482));
    ClkMux I__11777 (
            .O(N__49846),
            .I(N__49482));
    ClkMux I__11776 (
            .O(N__49845),
            .I(N__49482));
    ClkMux I__11775 (
            .O(N__49844),
            .I(N__49482));
    ClkMux I__11774 (
            .O(N__49843),
            .I(N__49482));
    ClkMux I__11773 (
            .O(N__49842),
            .I(N__49482));
    ClkMux I__11772 (
            .O(N__49841),
            .I(N__49482));
    ClkMux I__11771 (
            .O(N__49840),
            .I(N__49482));
    ClkMux I__11770 (
            .O(N__49839),
            .I(N__49482));
    ClkMux I__11769 (
            .O(N__49838),
            .I(N__49482));
    ClkMux I__11768 (
            .O(N__49837),
            .I(N__49482));
    ClkMux I__11767 (
            .O(N__49836),
            .I(N__49482));
    ClkMux I__11766 (
            .O(N__49835),
            .I(N__49482));
    ClkMux I__11765 (
            .O(N__49834),
            .I(N__49482));
    ClkMux I__11764 (
            .O(N__49833),
            .I(N__49482));
    ClkMux I__11763 (
            .O(N__49832),
            .I(N__49482));
    ClkMux I__11762 (
            .O(N__49831),
            .I(N__49482));
    ClkMux I__11761 (
            .O(N__49830),
            .I(N__49482));
    ClkMux I__11760 (
            .O(N__49829),
            .I(N__49482));
    ClkMux I__11759 (
            .O(N__49828),
            .I(N__49482));
    ClkMux I__11758 (
            .O(N__49827),
            .I(N__49482));
    ClkMux I__11757 (
            .O(N__49826),
            .I(N__49482));
    ClkMux I__11756 (
            .O(N__49825),
            .I(N__49482));
    ClkMux I__11755 (
            .O(N__49824),
            .I(N__49482));
    ClkMux I__11754 (
            .O(N__49823),
            .I(N__49482));
    ClkMux I__11753 (
            .O(N__49822),
            .I(N__49482));
    ClkMux I__11752 (
            .O(N__49821),
            .I(N__49482));
    ClkMux I__11751 (
            .O(N__49820),
            .I(N__49482));
    ClkMux I__11750 (
            .O(N__49819),
            .I(N__49482));
    ClkMux I__11749 (
            .O(N__49818),
            .I(N__49482));
    ClkMux I__11748 (
            .O(N__49817),
            .I(N__49482));
    ClkMux I__11747 (
            .O(N__49816),
            .I(N__49482));
    ClkMux I__11746 (
            .O(N__49815),
            .I(N__49482));
    ClkMux I__11745 (
            .O(N__49814),
            .I(N__49482));
    ClkMux I__11744 (
            .O(N__49813),
            .I(N__49482));
    ClkMux I__11743 (
            .O(N__49812),
            .I(N__49482));
    ClkMux I__11742 (
            .O(N__49811),
            .I(N__49482));
    ClkMux I__11741 (
            .O(N__49810),
            .I(N__49482));
    ClkMux I__11740 (
            .O(N__49809),
            .I(N__49482));
    ClkMux I__11739 (
            .O(N__49808),
            .I(N__49482));
    ClkMux I__11738 (
            .O(N__49807),
            .I(N__49482));
    ClkMux I__11737 (
            .O(N__49806),
            .I(N__49482));
    ClkMux I__11736 (
            .O(N__49805),
            .I(N__49482));
    ClkMux I__11735 (
            .O(N__49804),
            .I(N__49482));
    ClkMux I__11734 (
            .O(N__49803),
            .I(N__49482));
    ClkMux I__11733 (
            .O(N__49802),
            .I(N__49482));
    ClkMux I__11732 (
            .O(N__49801),
            .I(N__49482));
    ClkMux I__11731 (
            .O(N__49800),
            .I(N__49482));
    ClkMux I__11730 (
            .O(N__49799),
            .I(N__49482));
    GlobalMux I__11729 (
            .O(N__49482),
            .I(clk_100mhz_0));
    InMux I__11728 (
            .O(N__49479),
            .I(N__49473));
    InMux I__11727 (
            .O(N__49478),
            .I(N__49470));
    InMux I__11726 (
            .O(N__49477),
            .I(N__49467));
    InMux I__11725 (
            .O(N__49476),
            .I(N__49464));
    LocalMux I__11724 (
            .O(N__49473),
            .I(N__49461));
    LocalMux I__11723 (
            .O(N__49470),
            .I(N__49458));
    LocalMux I__11722 (
            .O(N__49467),
            .I(N__49455));
    LocalMux I__11721 (
            .O(N__49464),
            .I(N__49447));
    Glb2LocalMux I__11720 (
            .O(N__49461),
            .I(N__48960));
    Glb2LocalMux I__11719 (
            .O(N__49458),
            .I(N__48960));
    Glb2LocalMux I__11718 (
            .O(N__49455),
            .I(N__48960));
    SRMux I__11717 (
            .O(N__49454),
            .I(N__48960));
    SRMux I__11716 (
            .O(N__49453),
            .I(N__48960));
    SRMux I__11715 (
            .O(N__49452),
            .I(N__48960));
    SRMux I__11714 (
            .O(N__49451),
            .I(N__48960));
    SRMux I__11713 (
            .O(N__49450),
            .I(N__48960));
    Glb2LocalMux I__11712 (
            .O(N__49447),
            .I(N__48960));
    SRMux I__11711 (
            .O(N__49446),
            .I(N__48960));
    SRMux I__11710 (
            .O(N__49445),
            .I(N__48960));
    SRMux I__11709 (
            .O(N__49444),
            .I(N__48960));
    SRMux I__11708 (
            .O(N__49443),
            .I(N__48960));
    SRMux I__11707 (
            .O(N__49442),
            .I(N__48960));
    SRMux I__11706 (
            .O(N__49441),
            .I(N__48960));
    SRMux I__11705 (
            .O(N__49440),
            .I(N__48960));
    SRMux I__11704 (
            .O(N__49439),
            .I(N__48960));
    SRMux I__11703 (
            .O(N__49438),
            .I(N__48960));
    SRMux I__11702 (
            .O(N__49437),
            .I(N__48960));
    SRMux I__11701 (
            .O(N__49436),
            .I(N__48960));
    SRMux I__11700 (
            .O(N__49435),
            .I(N__48960));
    SRMux I__11699 (
            .O(N__49434),
            .I(N__48960));
    SRMux I__11698 (
            .O(N__49433),
            .I(N__48960));
    SRMux I__11697 (
            .O(N__49432),
            .I(N__48960));
    SRMux I__11696 (
            .O(N__49431),
            .I(N__48960));
    SRMux I__11695 (
            .O(N__49430),
            .I(N__48960));
    SRMux I__11694 (
            .O(N__49429),
            .I(N__48960));
    SRMux I__11693 (
            .O(N__49428),
            .I(N__48960));
    SRMux I__11692 (
            .O(N__49427),
            .I(N__48960));
    SRMux I__11691 (
            .O(N__49426),
            .I(N__48960));
    SRMux I__11690 (
            .O(N__49425),
            .I(N__48960));
    SRMux I__11689 (
            .O(N__49424),
            .I(N__48960));
    SRMux I__11688 (
            .O(N__49423),
            .I(N__48960));
    SRMux I__11687 (
            .O(N__49422),
            .I(N__48960));
    SRMux I__11686 (
            .O(N__49421),
            .I(N__48960));
    SRMux I__11685 (
            .O(N__49420),
            .I(N__48960));
    SRMux I__11684 (
            .O(N__49419),
            .I(N__48960));
    SRMux I__11683 (
            .O(N__49418),
            .I(N__48960));
    SRMux I__11682 (
            .O(N__49417),
            .I(N__48960));
    SRMux I__11681 (
            .O(N__49416),
            .I(N__48960));
    SRMux I__11680 (
            .O(N__49415),
            .I(N__48960));
    SRMux I__11679 (
            .O(N__49414),
            .I(N__48960));
    SRMux I__11678 (
            .O(N__49413),
            .I(N__48960));
    SRMux I__11677 (
            .O(N__49412),
            .I(N__48960));
    SRMux I__11676 (
            .O(N__49411),
            .I(N__48960));
    SRMux I__11675 (
            .O(N__49410),
            .I(N__48960));
    SRMux I__11674 (
            .O(N__49409),
            .I(N__48960));
    SRMux I__11673 (
            .O(N__49408),
            .I(N__48960));
    SRMux I__11672 (
            .O(N__49407),
            .I(N__48960));
    SRMux I__11671 (
            .O(N__49406),
            .I(N__48960));
    SRMux I__11670 (
            .O(N__49405),
            .I(N__48960));
    SRMux I__11669 (
            .O(N__49404),
            .I(N__48960));
    SRMux I__11668 (
            .O(N__49403),
            .I(N__48960));
    SRMux I__11667 (
            .O(N__49402),
            .I(N__48960));
    SRMux I__11666 (
            .O(N__49401),
            .I(N__48960));
    SRMux I__11665 (
            .O(N__49400),
            .I(N__48960));
    SRMux I__11664 (
            .O(N__49399),
            .I(N__48960));
    SRMux I__11663 (
            .O(N__49398),
            .I(N__48960));
    SRMux I__11662 (
            .O(N__49397),
            .I(N__48960));
    SRMux I__11661 (
            .O(N__49396),
            .I(N__48960));
    SRMux I__11660 (
            .O(N__49395),
            .I(N__48960));
    SRMux I__11659 (
            .O(N__49394),
            .I(N__48960));
    SRMux I__11658 (
            .O(N__49393),
            .I(N__48960));
    SRMux I__11657 (
            .O(N__49392),
            .I(N__48960));
    SRMux I__11656 (
            .O(N__49391),
            .I(N__48960));
    SRMux I__11655 (
            .O(N__49390),
            .I(N__48960));
    SRMux I__11654 (
            .O(N__49389),
            .I(N__48960));
    SRMux I__11653 (
            .O(N__49388),
            .I(N__48960));
    SRMux I__11652 (
            .O(N__49387),
            .I(N__48960));
    SRMux I__11651 (
            .O(N__49386),
            .I(N__48960));
    SRMux I__11650 (
            .O(N__49385),
            .I(N__48960));
    SRMux I__11649 (
            .O(N__49384),
            .I(N__48960));
    SRMux I__11648 (
            .O(N__49383),
            .I(N__48960));
    SRMux I__11647 (
            .O(N__49382),
            .I(N__48960));
    SRMux I__11646 (
            .O(N__49381),
            .I(N__48960));
    SRMux I__11645 (
            .O(N__49380),
            .I(N__48960));
    SRMux I__11644 (
            .O(N__49379),
            .I(N__48960));
    SRMux I__11643 (
            .O(N__49378),
            .I(N__48960));
    SRMux I__11642 (
            .O(N__49377),
            .I(N__48960));
    SRMux I__11641 (
            .O(N__49376),
            .I(N__48960));
    SRMux I__11640 (
            .O(N__49375),
            .I(N__48960));
    SRMux I__11639 (
            .O(N__49374),
            .I(N__48960));
    SRMux I__11638 (
            .O(N__49373),
            .I(N__48960));
    SRMux I__11637 (
            .O(N__49372),
            .I(N__48960));
    SRMux I__11636 (
            .O(N__49371),
            .I(N__48960));
    SRMux I__11635 (
            .O(N__49370),
            .I(N__48960));
    SRMux I__11634 (
            .O(N__49369),
            .I(N__48960));
    SRMux I__11633 (
            .O(N__49368),
            .I(N__48960));
    SRMux I__11632 (
            .O(N__49367),
            .I(N__48960));
    SRMux I__11631 (
            .O(N__49366),
            .I(N__48960));
    SRMux I__11630 (
            .O(N__49365),
            .I(N__48960));
    SRMux I__11629 (
            .O(N__49364),
            .I(N__48960));
    SRMux I__11628 (
            .O(N__49363),
            .I(N__48960));
    SRMux I__11627 (
            .O(N__49362),
            .I(N__48960));
    SRMux I__11626 (
            .O(N__49361),
            .I(N__48960));
    SRMux I__11625 (
            .O(N__49360),
            .I(N__48960));
    SRMux I__11624 (
            .O(N__49359),
            .I(N__48960));
    SRMux I__11623 (
            .O(N__49358),
            .I(N__48960));
    SRMux I__11622 (
            .O(N__49357),
            .I(N__48960));
    SRMux I__11621 (
            .O(N__49356),
            .I(N__48960));
    SRMux I__11620 (
            .O(N__49355),
            .I(N__48960));
    SRMux I__11619 (
            .O(N__49354),
            .I(N__48960));
    SRMux I__11618 (
            .O(N__49353),
            .I(N__48960));
    SRMux I__11617 (
            .O(N__49352),
            .I(N__48960));
    SRMux I__11616 (
            .O(N__49351),
            .I(N__48960));
    SRMux I__11615 (
            .O(N__49350),
            .I(N__48960));
    SRMux I__11614 (
            .O(N__49349),
            .I(N__48960));
    SRMux I__11613 (
            .O(N__49348),
            .I(N__48960));
    SRMux I__11612 (
            .O(N__49347),
            .I(N__48960));
    SRMux I__11611 (
            .O(N__49346),
            .I(N__48960));
    SRMux I__11610 (
            .O(N__49345),
            .I(N__48960));
    SRMux I__11609 (
            .O(N__49344),
            .I(N__48960));
    SRMux I__11608 (
            .O(N__49343),
            .I(N__48960));
    SRMux I__11607 (
            .O(N__49342),
            .I(N__48960));
    SRMux I__11606 (
            .O(N__49341),
            .I(N__48960));
    SRMux I__11605 (
            .O(N__49340),
            .I(N__48960));
    SRMux I__11604 (
            .O(N__49339),
            .I(N__48960));
    SRMux I__11603 (
            .O(N__49338),
            .I(N__48960));
    SRMux I__11602 (
            .O(N__49337),
            .I(N__48960));
    SRMux I__11601 (
            .O(N__49336),
            .I(N__48960));
    SRMux I__11600 (
            .O(N__49335),
            .I(N__48960));
    SRMux I__11599 (
            .O(N__49334),
            .I(N__48960));
    SRMux I__11598 (
            .O(N__49333),
            .I(N__48960));
    SRMux I__11597 (
            .O(N__49332),
            .I(N__48960));
    SRMux I__11596 (
            .O(N__49331),
            .I(N__48960));
    SRMux I__11595 (
            .O(N__49330),
            .I(N__48960));
    SRMux I__11594 (
            .O(N__49329),
            .I(N__48960));
    SRMux I__11593 (
            .O(N__49328),
            .I(N__48960));
    SRMux I__11592 (
            .O(N__49327),
            .I(N__48960));
    SRMux I__11591 (
            .O(N__49326),
            .I(N__48960));
    SRMux I__11590 (
            .O(N__49325),
            .I(N__48960));
    SRMux I__11589 (
            .O(N__49324),
            .I(N__48960));
    SRMux I__11588 (
            .O(N__49323),
            .I(N__48960));
    SRMux I__11587 (
            .O(N__49322),
            .I(N__48960));
    SRMux I__11586 (
            .O(N__49321),
            .I(N__48960));
    SRMux I__11585 (
            .O(N__49320),
            .I(N__48960));
    SRMux I__11584 (
            .O(N__49319),
            .I(N__48960));
    SRMux I__11583 (
            .O(N__49318),
            .I(N__48960));
    SRMux I__11582 (
            .O(N__49317),
            .I(N__48960));
    SRMux I__11581 (
            .O(N__49316),
            .I(N__48960));
    SRMux I__11580 (
            .O(N__49315),
            .I(N__48960));
    SRMux I__11579 (
            .O(N__49314),
            .I(N__48960));
    SRMux I__11578 (
            .O(N__49313),
            .I(N__48960));
    SRMux I__11577 (
            .O(N__49312),
            .I(N__48960));
    SRMux I__11576 (
            .O(N__49311),
            .I(N__48960));
    SRMux I__11575 (
            .O(N__49310),
            .I(N__48960));
    SRMux I__11574 (
            .O(N__49309),
            .I(N__48960));
    SRMux I__11573 (
            .O(N__49308),
            .I(N__48960));
    SRMux I__11572 (
            .O(N__49307),
            .I(N__48960));
    SRMux I__11571 (
            .O(N__49306),
            .I(N__48960));
    SRMux I__11570 (
            .O(N__49305),
            .I(N__48960));
    SRMux I__11569 (
            .O(N__49304),
            .I(N__48960));
    SRMux I__11568 (
            .O(N__49303),
            .I(N__48960));
    SRMux I__11567 (
            .O(N__49302),
            .I(N__48960));
    SRMux I__11566 (
            .O(N__49301),
            .I(N__48960));
    SRMux I__11565 (
            .O(N__49300),
            .I(N__48960));
    SRMux I__11564 (
            .O(N__49299),
            .I(N__48960));
    SRMux I__11563 (
            .O(N__49298),
            .I(N__48960));
    SRMux I__11562 (
            .O(N__49297),
            .I(N__48960));
    SRMux I__11561 (
            .O(N__49296),
            .I(N__48960));
    SRMux I__11560 (
            .O(N__49295),
            .I(N__48960));
    SRMux I__11559 (
            .O(N__49294),
            .I(N__48960));
    SRMux I__11558 (
            .O(N__49293),
            .I(N__48960));
    SRMux I__11557 (
            .O(N__49292),
            .I(N__48960));
    SRMux I__11556 (
            .O(N__49291),
            .I(N__48960));
    GlobalMux I__11555 (
            .O(N__48960),
            .I(N__48957));
    gio2CtrlBuf I__11554 (
            .O(N__48957),
            .I(red_c_g));
    InMux I__11553 (
            .O(N__48954),
            .I(N__48948));
    CascadeMux I__11552 (
            .O(N__48953),
            .I(N__48945));
    CascadeMux I__11551 (
            .O(N__48952),
            .I(N__48941));
    CascadeMux I__11550 (
            .O(N__48951),
            .I(N__48937));
    LocalMux I__11549 (
            .O(N__48948),
            .I(N__48933));
    InMux I__11548 (
            .O(N__48945),
            .I(N__48919));
    InMux I__11547 (
            .O(N__48944),
            .I(N__48919));
    InMux I__11546 (
            .O(N__48941),
            .I(N__48919));
    InMux I__11545 (
            .O(N__48940),
            .I(N__48919));
    InMux I__11544 (
            .O(N__48937),
            .I(N__48919));
    InMux I__11543 (
            .O(N__48936),
            .I(N__48919));
    Span12Mux_s7_v I__11542 (
            .O(N__48933),
            .I(N__48916));
    InMux I__11541 (
            .O(N__48932),
            .I(N__48913));
    LocalMux I__11540 (
            .O(N__48919),
            .I(N__48910));
    Span12Mux_h I__11539 (
            .O(N__48916),
            .I(N__48905));
    LocalMux I__11538 (
            .O(N__48913),
            .I(N__48905));
    Span4Mux_h I__11537 (
            .O(N__48910),
            .I(N__48902));
    Span12Mux_h I__11536 (
            .O(N__48905),
            .I(N__48899));
    Span4Mux_h I__11535 (
            .O(N__48902),
            .I(N__48896));
    Odrv12 I__11534 (
            .O(N__48899),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    Odrv4 I__11533 (
            .O(N__48896),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    InMux I__11532 (
            .O(N__48891),
            .I(N__48888));
    LocalMux I__11531 (
            .O(N__48888),
            .I(N__48885));
    Span12Mux_v I__11530 (
            .O(N__48885),
            .I(N__48882));
    Span12Mux_h I__11529 (
            .O(N__48882),
            .I(N__48878));
    InMux I__11528 (
            .O(N__48881),
            .I(N__48875));
    Odrv12 I__11527 (
            .O(N__48878),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    LocalMux I__11526 (
            .O(N__48875),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    CascadeMux I__11525 (
            .O(N__48870),
            .I(N__48846));
    CascadeMux I__11524 (
            .O(N__48869),
            .I(N__48843));
    InMux I__11523 (
            .O(N__48868),
            .I(N__48840));
    InMux I__11522 (
            .O(N__48867),
            .I(N__48818));
    InMux I__11521 (
            .O(N__48866),
            .I(N__48818));
    InMux I__11520 (
            .O(N__48865),
            .I(N__48818));
    InMux I__11519 (
            .O(N__48864),
            .I(N__48818));
    InMux I__11518 (
            .O(N__48863),
            .I(N__48818));
    InMux I__11517 (
            .O(N__48862),
            .I(N__48818));
    InMux I__11516 (
            .O(N__48861),
            .I(N__48818));
    InMux I__11515 (
            .O(N__48860),
            .I(N__48818));
    InMux I__11514 (
            .O(N__48859),
            .I(N__48803));
    InMux I__11513 (
            .O(N__48858),
            .I(N__48803));
    InMux I__11512 (
            .O(N__48857),
            .I(N__48803));
    InMux I__11511 (
            .O(N__48856),
            .I(N__48803));
    InMux I__11510 (
            .O(N__48855),
            .I(N__48803));
    InMux I__11509 (
            .O(N__48854),
            .I(N__48803));
    InMux I__11508 (
            .O(N__48853),
            .I(N__48803));
    CascadeMux I__11507 (
            .O(N__48852),
            .I(N__48800));
    CascadeMux I__11506 (
            .O(N__48851),
            .I(N__48797));
    CascadeMux I__11505 (
            .O(N__48850),
            .I(N__48793));
    CascadeMux I__11504 (
            .O(N__48849),
            .I(N__48790));
    InMux I__11503 (
            .O(N__48846),
            .I(N__48785));
    InMux I__11502 (
            .O(N__48843),
            .I(N__48785));
    LocalMux I__11501 (
            .O(N__48840),
            .I(N__48782));
    InMux I__11500 (
            .O(N__48839),
            .I(N__48775));
    InMux I__11499 (
            .O(N__48838),
            .I(N__48775));
    InMux I__11498 (
            .O(N__48837),
            .I(N__48768));
    InMux I__11497 (
            .O(N__48836),
            .I(N__48768));
    InMux I__11496 (
            .O(N__48835),
            .I(N__48768));
    LocalMux I__11495 (
            .O(N__48818),
            .I(N__48763));
    LocalMux I__11494 (
            .O(N__48803),
            .I(N__48763));
    InMux I__11493 (
            .O(N__48800),
            .I(N__48758));
    InMux I__11492 (
            .O(N__48797),
            .I(N__48758));
    InMux I__11491 (
            .O(N__48796),
            .I(N__48751));
    InMux I__11490 (
            .O(N__48793),
            .I(N__48751));
    InMux I__11489 (
            .O(N__48790),
            .I(N__48751));
    LocalMux I__11488 (
            .O(N__48785),
            .I(N__48748));
    Span4Mux_s3_h I__11487 (
            .O(N__48782),
            .I(N__48745));
    CascadeMux I__11486 (
            .O(N__48781),
            .I(N__48742));
    InMux I__11485 (
            .O(N__48780),
            .I(N__48739));
    LocalMux I__11484 (
            .O(N__48775),
            .I(N__48734));
    LocalMux I__11483 (
            .O(N__48768),
            .I(N__48734));
    Span4Mux_s3_h I__11482 (
            .O(N__48763),
            .I(N__48731));
    LocalMux I__11481 (
            .O(N__48758),
            .I(N__48722));
    LocalMux I__11480 (
            .O(N__48751),
            .I(N__48722));
    Span4Mux_h I__11479 (
            .O(N__48748),
            .I(N__48722));
    Span4Mux_h I__11478 (
            .O(N__48745),
            .I(N__48719));
    InMux I__11477 (
            .O(N__48742),
            .I(N__48716));
    LocalMux I__11476 (
            .O(N__48739),
            .I(N__48713));
    Span4Mux_s2_h I__11475 (
            .O(N__48734),
            .I(N__48710));
    Span4Mux_h I__11474 (
            .O(N__48731),
            .I(N__48707));
    CascadeMux I__11473 (
            .O(N__48730),
            .I(N__48704));
    CascadeMux I__11472 (
            .O(N__48729),
            .I(N__48701));
    Span4Mux_h I__11471 (
            .O(N__48722),
            .I(N__48696));
    Span4Mux_h I__11470 (
            .O(N__48719),
            .I(N__48696));
    LocalMux I__11469 (
            .O(N__48716),
            .I(N__48689));
    Span4Mux_h I__11468 (
            .O(N__48713),
            .I(N__48689));
    Span4Mux_h I__11467 (
            .O(N__48710),
            .I(N__48689));
    Span4Mux_h I__11466 (
            .O(N__48707),
            .I(N__48686));
    InMux I__11465 (
            .O(N__48704),
            .I(N__48683));
    InMux I__11464 (
            .O(N__48701),
            .I(N__48680));
    Span4Mux_h I__11463 (
            .O(N__48696),
            .I(N__48677));
    Span4Mux_h I__11462 (
            .O(N__48689),
            .I(N__48672));
    Span4Mux_h I__11461 (
            .O(N__48686),
            .I(N__48672));
    LocalMux I__11460 (
            .O(N__48683),
            .I(N_19_1));
    LocalMux I__11459 (
            .O(N__48680),
            .I(N_19_1));
    Odrv4 I__11458 (
            .O(N__48677),
            .I(N_19_1));
    Odrv4 I__11457 (
            .O(N__48672),
            .I(N_19_1));
    InMux I__11456 (
            .O(N__48663),
            .I(N__48660));
    LocalMux I__11455 (
            .O(N__48660),
            .I(N__48657));
    Span12Mux_s8_h I__11454 (
            .O(N__48657),
            .I(N__48654));
    Span12Mux_h I__11453 (
            .O(N__48654),
            .I(N__48651));
    Odrv12 I__11452 (
            .O(N__48651),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__11451 (
            .O(N__48648),
            .I(N__48629));
    InMux I__11450 (
            .O(N__48647),
            .I(N__48629));
    InMux I__11449 (
            .O(N__48646),
            .I(N__48629));
    InMux I__11448 (
            .O(N__48645),
            .I(N__48629));
    InMux I__11447 (
            .O(N__48644),
            .I(N__48619));
    InMux I__11446 (
            .O(N__48643),
            .I(N__48612));
    InMux I__11445 (
            .O(N__48642),
            .I(N__48612));
    InMux I__11444 (
            .O(N__48641),
            .I(N__48612));
    InMux I__11443 (
            .O(N__48640),
            .I(N__48607));
    InMux I__11442 (
            .O(N__48639),
            .I(N__48607));
    InMux I__11441 (
            .O(N__48638),
            .I(N__48604));
    LocalMux I__11440 (
            .O(N__48629),
            .I(N__48601));
    InMux I__11439 (
            .O(N__48628),
            .I(N__48592));
    InMux I__11438 (
            .O(N__48627),
            .I(N__48592));
    InMux I__11437 (
            .O(N__48626),
            .I(N__48592));
    InMux I__11436 (
            .O(N__48625),
            .I(N__48592));
    InMux I__11435 (
            .O(N__48624),
            .I(N__48585));
    InMux I__11434 (
            .O(N__48623),
            .I(N__48585));
    InMux I__11433 (
            .O(N__48622),
            .I(N__48585));
    LocalMux I__11432 (
            .O(N__48619),
            .I(N__48577));
    LocalMux I__11431 (
            .O(N__48612),
            .I(N__48574));
    LocalMux I__11430 (
            .O(N__48607),
            .I(N__48563));
    LocalMux I__11429 (
            .O(N__48604),
            .I(N__48563));
    Span4Mux_v I__11428 (
            .O(N__48601),
            .I(N__48563));
    LocalMux I__11427 (
            .O(N__48592),
            .I(N__48563));
    LocalMux I__11426 (
            .O(N__48585),
            .I(N__48563));
    InMux I__11425 (
            .O(N__48584),
            .I(N__48552));
    InMux I__11424 (
            .O(N__48583),
            .I(N__48552));
    InMux I__11423 (
            .O(N__48582),
            .I(N__48552));
    InMux I__11422 (
            .O(N__48581),
            .I(N__48552));
    InMux I__11421 (
            .O(N__48580),
            .I(N__48552));
    Span4Mux_h I__11420 (
            .O(N__48577),
            .I(N__48545));
    Span4Mux_v I__11419 (
            .O(N__48574),
            .I(N__48545));
    Span4Mux_v I__11418 (
            .O(N__48563),
            .I(N__48540));
    LocalMux I__11417 (
            .O(N__48552),
            .I(N__48540));
    InMux I__11416 (
            .O(N__48551),
            .I(N__48537));
    InMux I__11415 (
            .O(N__48550),
            .I(N__48534));
    Odrv4 I__11414 (
            .O(N__48545),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__11413 (
            .O(N__48540),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__11412 (
            .O(N__48537),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__11411 (
            .O(N__48534),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__11410 (
            .O(N__48525),
            .I(N__48520));
    InMux I__11409 (
            .O(N__48524),
            .I(N__48517));
    InMux I__11408 (
            .O(N__48523),
            .I(N__48514));
    LocalMux I__11407 (
            .O(N__48520),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__11406 (
            .O(N__48517),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__11405 (
            .O(N__48514),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__11404 (
            .O(N__48507),
            .I(N__48504));
    LocalMux I__11403 (
            .O(N__48504),
            .I(N__48498));
    InMux I__11402 (
            .O(N__48503),
            .I(N__48491));
    InMux I__11401 (
            .O(N__48502),
            .I(N__48491));
    InMux I__11400 (
            .O(N__48501),
            .I(N__48491));
    Odrv4 I__11399 (
            .O(N__48498),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__11398 (
            .O(N__48491),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__11397 (
            .O(N__48486),
            .I(N__48483));
    InMux I__11396 (
            .O(N__48483),
            .I(N__48480));
    LocalMux I__11395 (
            .O(N__48480),
            .I(N__48477));
    Span4Mux_v I__11394 (
            .O(N__48477),
            .I(N__48474));
    Span4Mux_h I__11393 (
            .O(N__48474),
            .I(N__48471));
    Odrv4 I__11392 (
            .O(N__48471),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__11391 (
            .O(N__48468),
            .I(N__48464));
    InMux I__11390 (
            .O(N__48467),
            .I(N__48461));
    LocalMux I__11389 (
            .O(N__48464),
            .I(N__48457));
    LocalMux I__11388 (
            .O(N__48461),
            .I(N__48454));
    InMux I__11387 (
            .O(N__48460),
            .I(N__48451));
    Span4Mux_h I__11386 (
            .O(N__48457),
            .I(N__48447));
    Span4Mux_v I__11385 (
            .O(N__48454),
            .I(N__48442));
    LocalMux I__11384 (
            .O(N__48451),
            .I(N__48442));
    InMux I__11383 (
            .O(N__48450),
            .I(N__48439));
    Odrv4 I__11382 (
            .O(N__48447),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__11381 (
            .O(N__48442),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__11380 (
            .O(N__48439),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    CascadeMux I__11379 (
            .O(N__48432),
            .I(N__48429));
    InMux I__11378 (
            .O(N__48429),
            .I(N__48426));
    LocalMux I__11377 (
            .O(N__48426),
            .I(N__48422));
    InMux I__11376 (
            .O(N__48425),
            .I(N__48418));
    Span4Mux_v I__11375 (
            .O(N__48422),
            .I(N__48415));
    InMux I__11374 (
            .O(N__48421),
            .I(N__48412));
    LocalMux I__11373 (
            .O(N__48418),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__11372 (
            .O(N__48415),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__11371 (
            .O(N__48412),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__11370 (
            .O(N__48405),
            .I(N__48402));
    InMux I__11369 (
            .O(N__48402),
            .I(N__48399));
    LocalMux I__11368 (
            .O(N__48399),
            .I(N__48396));
    Odrv12 I__11367 (
            .O(N__48396),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    InMux I__11366 (
            .O(N__48393),
            .I(N__48389));
    InMux I__11365 (
            .O(N__48392),
            .I(N__48386));
    LocalMux I__11364 (
            .O(N__48389),
            .I(N__48381));
    LocalMux I__11363 (
            .O(N__48386),
            .I(N__48378));
    InMux I__11362 (
            .O(N__48385),
            .I(N__48373));
    InMux I__11361 (
            .O(N__48384),
            .I(N__48373));
    Span4Mux_v I__11360 (
            .O(N__48381),
            .I(N__48368));
    Span4Mux_h I__11359 (
            .O(N__48378),
            .I(N__48368));
    LocalMux I__11358 (
            .O(N__48373),
            .I(N__48365));
    Odrv4 I__11357 (
            .O(N__48368),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__11356 (
            .O(N__48365),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__11355 (
            .O(N__48360),
            .I(N__48357));
    LocalMux I__11354 (
            .O(N__48357),
            .I(N__48354));
    Span4Mux_h I__11353 (
            .O(N__48354),
            .I(N__48349));
    InMux I__11352 (
            .O(N__48353),
            .I(N__48346));
    InMux I__11351 (
            .O(N__48352),
            .I(N__48343));
    Odrv4 I__11350 (
            .O(N__48349),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__11349 (
            .O(N__48346),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__11348 (
            .O(N__48343),
            .I(\current_shift_inst.un4_control_input1_11 ));
    CascadeMux I__11347 (
            .O(N__48336),
            .I(N__48333));
    InMux I__11346 (
            .O(N__48333),
            .I(N__48330));
    LocalMux I__11345 (
            .O(N__48330),
            .I(N__48327));
    Span4Mux_h I__11344 (
            .O(N__48327),
            .I(N__48324));
    Odrv4 I__11343 (
            .O(N__48324),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    CascadeMux I__11342 (
            .O(N__48321),
            .I(N__48318));
    InMux I__11341 (
            .O(N__48318),
            .I(N__48315));
    LocalMux I__11340 (
            .O(N__48315),
            .I(N__48310));
    InMux I__11339 (
            .O(N__48314),
            .I(N__48305));
    InMux I__11338 (
            .O(N__48313),
            .I(N__48305));
    Span4Mux_h I__11337 (
            .O(N__48310),
            .I(N__48299));
    LocalMux I__11336 (
            .O(N__48305),
            .I(N__48299));
    InMux I__11335 (
            .O(N__48304),
            .I(N__48296));
    Odrv4 I__11334 (
            .O(N__48299),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__11333 (
            .O(N__48296),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    CascadeMux I__11332 (
            .O(N__48291),
            .I(N__48288));
    InMux I__11331 (
            .O(N__48288),
            .I(N__48283));
    InMux I__11330 (
            .O(N__48287),
            .I(N__48280));
    InMux I__11329 (
            .O(N__48286),
            .I(N__48277));
    LocalMux I__11328 (
            .O(N__48283),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__11327 (
            .O(N__48280),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__11326 (
            .O(N__48277),
            .I(\current_shift_inst.un4_control_input1_21 ));
    CascadeMux I__11325 (
            .O(N__48270),
            .I(N__48267));
    InMux I__11324 (
            .O(N__48267),
            .I(N__48264));
    LocalMux I__11323 (
            .O(N__48264),
            .I(N__48261));
    Span4Mux_h I__11322 (
            .O(N__48261),
            .I(N__48258));
    Odrv4 I__11321 (
            .O(N__48258),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__11320 (
            .O(N__48255),
            .I(N__48248));
    InMux I__11319 (
            .O(N__48254),
            .I(N__48245));
    InMux I__11318 (
            .O(N__48253),
            .I(N__48229));
    InMux I__11317 (
            .O(N__48252),
            .I(N__48229));
    CascadeMux I__11316 (
            .O(N__48251),
            .I(N__48217));
    LocalMux I__11315 (
            .O(N__48248),
            .I(N__48202));
    LocalMux I__11314 (
            .O(N__48245),
            .I(N__48199));
    InMux I__11313 (
            .O(N__48244),
            .I(N__48191));
    InMux I__11312 (
            .O(N__48243),
            .I(N__48191));
    InMux I__11311 (
            .O(N__48242),
            .I(N__48188));
    InMux I__11310 (
            .O(N__48241),
            .I(N__48170));
    InMux I__11309 (
            .O(N__48240),
            .I(N__48170));
    InMux I__11308 (
            .O(N__48239),
            .I(N__48170));
    InMux I__11307 (
            .O(N__48238),
            .I(N__48170));
    InMux I__11306 (
            .O(N__48237),
            .I(N__48159));
    InMux I__11305 (
            .O(N__48236),
            .I(N__48159));
    InMux I__11304 (
            .O(N__48235),
            .I(N__48154));
    InMux I__11303 (
            .O(N__48234),
            .I(N__48154));
    LocalMux I__11302 (
            .O(N__48229),
            .I(N__48151));
    InMux I__11301 (
            .O(N__48228),
            .I(N__48142));
    InMux I__11300 (
            .O(N__48227),
            .I(N__48142));
    InMux I__11299 (
            .O(N__48226),
            .I(N__48142));
    InMux I__11298 (
            .O(N__48225),
            .I(N__48142));
    InMux I__11297 (
            .O(N__48224),
            .I(N__48127));
    InMux I__11296 (
            .O(N__48223),
            .I(N__48127));
    InMux I__11295 (
            .O(N__48222),
            .I(N__48127));
    InMux I__11294 (
            .O(N__48221),
            .I(N__48127));
    InMux I__11293 (
            .O(N__48220),
            .I(N__48127));
    InMux I__11292 (
            .O(N__48217),
            .I(N__48127));
    InMux I__11291 (
            .O(N__48216),
            .I(N__48127));
    InMux I__11290 (
            .O(N__48215),
            .I(N__48110));
    InMux I__11289 (
            .O(N__48214),
            .I(N__48110));
    InMux I__11288 (
            .O(N__48213),
            .I(N__48110));
    InMux I__11287 (
            .O(N__48212),
            .I(N__48110));
    InMux I__11286 (
            .O(N__48211),
            .I(N__48110));
    InMux I__11285 (
            .O(N__48210),
            .I(N__48110));
    InMux I__11284 (
            .O(N__48209),
            .I(N__48110));
    InMux I__11283 (
            .O(N__48208),
            .I(N__48110));
    InMux I__11282 (
            .O(N__48207),
            .I(N__48107));
    InMux I__11281 (
            .O(N__48206),
            .I(N__48104));
    InMux I__11280 (
            .O(N__48205),
            .I(N__48101));
    Span4Mux_v I__11279 (
            .O(N__48202),
            .I(N__48098));
    Span4Mux_v I__11278 (
            .O(N__48199),
            .I(N__48095));
    CascadeMux I__11277 (
            .O(N__48198),
            .I(N__48088));
    InMux I__11276 (
            .O(N__48197),
            .I(N__48074));
    InMux I__11275 (
            .O(N__48196),
            .I(N__48074));
    LocalMux I__11274 (
            .O(N__48191),
            .I(N__48071));
    LocalMux I__11273 (
            .O(N__48188),
            .I(N__48068));
    InMux I__11272 (
            .O(N__48187),
            .I(N__48061));
    InMux I__11271 (
            .O(N__48186),
            .I(N__48061));
    InMux I__11270 (
            .O(N__48185),
            .I(N__48061));
    InMux I__11269 (
            .O(N__48184),
            .I(N__48056));
    InMux I__11268 (
            .O(N__48183),
            .I(N__48056));
    InMux I__11267 (
            .O(N__48182),
            .I(N__48047));
    InMux I__11266 (
            .O(N__48181),
            .I(N__48047));
    InMux I__11265 (
            .O(N__48180),
            .I(N__48047));
    InMux I__11264 (
            .O(N__48179),
            .I(N__48047));
    LocalMux I__11263 (
            .O(N__48170),
            .I(N__48044));
    InMux I__11262 (
            .O(N__48169),
            .I(N__48031));
    InMux I__11261 (
            .O(N__48168),
            .I(N__48031));
    InMux I__11260 (
            .O(N__48167),
            .I(N__48031));
    InMux I__11259 (
            .O(N__48166),
            .I(N__48031));
    InMux I__11258 (
            .O(N__48165),
            .I(N__48031));
    InMux I__11257 (
            .O(N__48164),
            .I(N__48031));
    LocalMux I__11256 (
            .O(N__48159),
            .I(N__48016));
    LocalMux I__11255 (
            .O(N__48154),
            .I(N__48016));
    Span4Mux_v I__11254 (
            .O(N__48151),
            .I(N__48016));
    LocalMux I__11253 (
            .O(N__48142),
            .I(N__48016));
    LocalMux I__11252 (
            .O(N__48127),
            .I(N__48016));
    LocalMux I__11251 (
            .O(N__48110),
            .I(N__48016));
    LocalMux I__11250 (
            .O(N__48107),
            .I(N__48016));
    LocalMux I__11249 (
            .O(N__48104),
            .I(N__48011));
    LocalMux I__11248 (
            .O(N__48101),
            .I(N__48011));
    Span4Mux_h I__11247 (
            .O(N__48098),
            .I(N__48003));
    Span4Mux_h I__11246 (
            .O(N__48095),
            .I(N__48003));
    InMux I__11245 (
            .O(N__48094),
            .I(N__47998));
    InMux I__11244 (
            .O(N__48093),
            .I(N__47998));
    InMux I__11243 (
            .O(N__48092),
            .I(N__47995));
    InMux I__11242 (
            .O(N__48091),
            .I(N__47990));
    InMux I__11241 (
            .O(N__48088),
            .I(N__47990));
    InMux I__11240 (
            .O(N__48087),
            .I(N__47987));
    InMux I__11239 (
            .O(N__48086),
            .I(N__47984));
    InMux I__11238 (
            .O(N__48085),
            .I(N__47969));
    InMux I__11237 (
            .O(N__48084),
            .I(N__47969));
    InMux I__11236 (
            .O(N__48083),
            .I(N__47969));
    InMux I__11235 (
            .O(N__48082),
            .I(N__47969));
    InMux I__11234 (
            .O(N__48081),
            .I(N__47969));
    InMux I__11233 (
            .O(N__48080),
            .I(N__47969));
    InMux I__11232 (
            .O(N__48079),
            .I(N__47969));
    LocalMux I__11231 (
            .O(N__48074),
            .I(N__47956));
    Sp12to4 I__11230 (
            .O(N__48071),
            .I(N__47956));
    Sp12to4 I__11229 (
            .O(N__48068),
            .I(N__47956));
    LocalMux I__11228 (
            .O(N__48061),
            .I(N__47956));
    LocalMux I__11227 (
            .O(N__48056),
            .I(N__47956));
    LocalMux I__11226 (
            .O(N__48047),
            .I(N__47956));
    Span4Mux_v I__11225 (
            .O(N__48044),
            .I(N__47947));
    LocalMux I__11224 (
            .O(N__48031),
            .I(N__47947));
    Span4Mux_v I__11223 (
            .O(N__48016),
            .I(N__47947));
    Span4Mux_v I__11222 (
            .O(N__48011),
            .I(N__47947));
    InMux I__11221 (
            .O(N__48010),
            .I(N__47940));
    InMux I__11220 (
            .O(N__48009),
            .I(N__47940));
    InMux I__11219 (
            .O(N__48008),
            .I(N__47940));
    Odrv4 I__11218 (
            .O(N__48003),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11217 (
            .O(N__47998),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11216 (
            .O(N__47995),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11215 (
            .O(N__47990),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11214 (
            .O(N__47987),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11213 (
            .O(N__47984),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11212 (
            .O(N__47969),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__11211 (
            .O(N__47956),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11210 (
            .O(N__47947),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11209 (
            .O(N__47940),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__11208 (
            .O(N__47919),
            .I(N__47915));
    CascadeMux I__11207 (
            .O(N__47918),
            .I(N__47912));
    LocalMux I__11206 (
            .O(N__47915),
            .I(N__47908));
    InMux I__11205 (
            .O(N__47912),
            .I(N__47905));
    InMux I__11204 (
            .O(N__47911),
            .I(N__47902));
    Span4Mux_h I__11203 (
            .O(N__47908),
            .I(N__47898));
    LocalMux I__11202 (
            .O(N__47905),
            .I(N__47895));
    LocalMux I__11201 (
            .O(N__47902),
            .I(N__47892));
    InMux I__11200 (
            .O(N__47901),
            .I(N__47889));
    Odrv4 I__11199 (
            .O(N__47898),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv12 I__11198 (
            .O(N__47895),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__11197 (
            .O(N__47892),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__11196 (
            .O(N__47889),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    CascadeMux I__11195 (
            .O(N__47880),
            .I(N__47867));
    CascadeMux I__11194 (
            .O(N__47879),
            .I(N__47858));
    CascadeMux I__11193 (
            .O(N__47878),
            .I(N__47854));
    CascadeMux I__11192 (
            .O(N__47877),
            .I(N__47850));
    CascadeMux I__11191 (
            .O(N__47876),
            .I(N__47843));
    CascadeMux I__11190 (
            .O(N__47875),
            .I(N__47840));
    CascadeMux I__11189 (
            .O(N__47874),
            .I(N__47831));
    CascadeMux I__11188 (
            .O(N__47873),
            .I(N__47827));
    CascadeMux I__11187 (
            .O(N__47872),
            .I(N__47823));
    InMux I__11186 (
            .O(N__47871),
            .I(N__47802));
    InMux I__11185 (
            .O(N__47870),
            .I(N__47802));
    InMux I__11184 (
            .O(N__47867),
            .I(N__47792));
    CascadeMux I__11183 (
            .O(N__47866),
            .I(N__47788));
    CascadeMux I__11182 (
            .O(N__47865),
            .I(N__47785));
    CascadeMux I__11181 (
            .O(N__47864),
            .I(N__47782));
    InMux I__11180 (
            .O(N__47863),
            .I(N__47769));
    InMux I__11179 (
            .O(N__47862),
            .I(N__47769));
    InMux I__11178 (
            .O(N__47861),
            .I(N__47769));
    InMux I__11177 (
            .O(N__47858),
            .I(N__47769));
    InMux I__11176 (
            .O(N__47857),
            .I(N__47769));
    InMux I__11175 (
            .O(N__47854),
            .I(N__47769));
    InMux I__11174 (
            .O(N__47853),
            .I(N__47763));
    InMux I__11173 (
            .O(N__47850),
            .I(N__47763));
    InMux I__11172 (
            .O(N__47849),
            .I(N__47758));
    InMux I__11171 (
            .O(N__47848),
            .I(N__47758));
    CascadeMux I__11170 (
            .O(N__47847),
            .I(N__47751));
    CascadeMux I__11169 (
            .O(N__47846),
            .I(N__47747));
    InMux I__11168 (
            .O(N__47843),
            .I(N__47736));
    InMux I__11167 (
            .O(N__47840),
            .I(N__47733));
    CascadeMux I__11166 (
            .O(N__47839),
            .I(N__47730));
    CascadeMux I__11165 (
            .O(N__47838),
            .I(N__47726));
    CascadeMux I__11164 (
            .O(N__47837),
            .I(N__47722));
    CascadeMux I__11163 (
            .O(N__47836),
            .I(N__47718));
    InMux I__11162 (
            .O(N__47835),
            .I(N__47701));
    InMux I__11161 (
            .O(N__47834),
            .I(N__47701));
    InMux I__11160 (
            .O(N__47831),
            .I(N__47701));
    InMux I__11159 (
            .O(N__47830),
            .I(N__47701));
    InMux I__11158 (
            .O(N__47827),
            .I(N__47701));
    InMux I__11157 (
            .O(N__47826),
            .I(N__47701));
    InMux I__11156 (
            .O(N__47823),
            .I(N__47701));
    InMux I__11155 (
            .O(N__47822),
            .I(N__47701));
    CascadeMux I__11154 (
            .O(N__47821),
            .I(N__47698));
    CascadeMux I__11153 (
            .O(N__47820),
            .I(N__47694));
    CascadeMux I__11152 (
            .O(N__47819),
            .I(N__47690));
    CascadeMux I__11151 (
            .O(N__47818),
            .I(N__47686));
    CascadeMux I__11150 (
            .O(N__47817),
            .I(N__47682));
    CascadeMux I__11149 (
            .O(N__47816),
            .I(N__47678));
    CascadeMux I__11148 (
            .O(N__47815),
            .I(N__47674));
    CascadeMux I__11147 (
            .O(N__47814),
            .I(N__47670));
    CascadeMux I__11146 (
            .O(N__47813),
            .I(N__47666));
    CascadeMux I__11145 (
            .O(N__47812),
            .I(N__47662));
    CascadeMux I__11144 (
            .O(N__47811),
            .I(N__47658));
    CascadeMux I__11143 (
            .O(N__47810),
            .I(N__47654));
    CascadeMux I__11142 (
            .O(N__47809),
            .I(N__47650));
    CascadeMux I__11141 (
            .O(N__47808),
            .I(N__47646));
    CascadeMux I__11140 (
            .O(N__47807),
            .I(N__47642));
    LocalMux I__11139 (
            .O(N__47802),
            .I(N__47638));
    InMux I__11138 (
            .O(N__47801),
            .I(N__47631));
    InMux I__11137 (
            .O(N__47800),
            .I(N__47631));
    InMux I__11136 (
            .O(N__47799),
            .I(N__47631));
    InMux I__11135 (
            .O(N__47798),
            .I(N__47624));
    InMux I__11134 (
            .O(N__47797),
            .I(N__47624));
    InMux I__11133 (
            .O(N__47796),
            .I(N__47624));
    CascadeMux I__11132 (
            .O(N__47795),
            .I(N__47620));
    LocalMux I__11131 (
            .O(N__47792),
            .I(N__47607));
    InMux I__11130 (
            .O(N__47791),
            .I(N__47604));
    InMux I__11129 (
            .O(N__47788),
            .I(N__47597));
    InMux I__11128 (
            .O(N__47785),
            .I(N__47597));
    InMux I__11127 (
            .O(N__47782),
            .I(N__47597));
    LocalMux I__11126 (
            .O(N__47769),
            .I(N__47594));
    InMux I__11125 (
            .O(N__47768),
            .I(N__47591));
    LocalMux I__11124 (
            .O(N__47763),
            .I(N__47579));
    LocalMux I__11123 (
            .O(N__47758),
            .I(N__47579));
    InMux I__11122 (
            .O(N__47757),
            .I(N__47564));
    InMux I__11121 (
            .O(N__47756),
            .I(N__47564));
    InMux I__11120 (
            .O(N__47755),
            .I(N__47564));
    InMux I__11119 (
            .O(N__47754),
            .I(N__47564));
    InMux I__11118 (
            .O(N__47751),
            .I(N__47564));
    InMux I__11117 (
            .O(N__47750),
            .I(N__47564));
    InMux I__11116 (
            .O(N__47747),
            .I(N__47564));
    InMux I__11115 (
            .O(N__47746),
            .I(N__47547));
    InMux I__11114 (
            .O(N__47745),
            .I(N__47547));
    InMux I__11113 (
            .O(N__47744),
            .I(N__47547));
    InMux I__11112 (
            .O(N__47743),
            .I(N__47547));
    InMux I__11111 (
            .O(N__47742),
            .I(N__47547));
    InMux I__11110 (
            .O(N__47741),
            .I(N__47547));
    InMux I__11109 (
            .O(N__47740),
            .I(N__47547));
    InMux I__11108 (
            .O(N__47739),
            .I(N__47547));
    LocalMux I__11107 (
            .O(N__47736),
            .I(N__47542));
    LocalMux I__11106 (
            .O(N__47733),
            .I(N__47542));
    InMux I__11105 (
            .O(N__47730),
            .I(N__47527));
    InMux I__11104 (
            .O(N__47729),
            .I(N__47527));
    InMux I__11103 (
            .O(N__47726),
            .I(N__47527));
    InMux I__11102 (
            .O(N__47725),
            .I(N__47527));
    InMux I__11101 (
            .O(N__47722),
            .I(N__47527));
    InMux I__11100 (
            .O(N__47721),
            .I(N__47527));
    InMux I__11099 (
            .O(N__47718),
            .I(N__47527));
    LocalMux I__11098 (
            .O(N__47701),
            .I(N__47524));
    InMux I__11097 (
            .O(N__47698),
            .I(N__47507));
    InMux I__11096 (
            .O(N__47697),
            .I(N__47507));
    InMux I__11095 (
            .O(N__47694),
            .I(N__47507));
    InMux I__11094 (
            .O(N__47693),
            .I(N__47507));
    InMux I__11093 (
            .O(N__47690),
            .I(N__47507));
    InMux I__11092 (
            .O(N__47689),
            .I(N__47507));
    InMux I__11091 (
            .O(N__47686),
            .I(N__47507));
    InMux I__11090 (
            .O(N__47685),
            .I(N__47507));
    InMux I__11089 (
            .O(N__47682),
            .I(N__47490));
    InMux I__11088 (
            .O(N__47681),
            .I(N__47490));
    InMux I__11087 (
            .O(N__47678),
            .I(N__47490));
    InMux I__11086 (
            .O(N__47677),
            .I(N__47490));
    InMux I__11085 (
            .O(N__47674),
            .I(N__47490));
    InMux I__11084 (
            .O(N__47673),
            .I(N__47490));
    InMux I__11083 (
            .O(N__47670),
            .I(N__47490));
    InMux I__11082 (
            .O(N__47669),
            .I(N__47490));
    InMux I__11081 (
            .O(N__47666),
            .I(N__47473));
    InMux I__11080 (
            .O(N__47665),
            .I(N__47473));
    InMux I__11079 (
            .O(N__47662),
            .I(N__47473));
    InMux I__11078 (
            .O(N__47661),
            .I(N__47473));
    InMux I__11077 (
            .O(N__47658),
            .I(N__47473));
    InMux I__11076 (
            .O(N__47657),
            .I(N__47473));
    InMux I__11075 (
            .O(N__47654),
            .I(N__47473));
    InMux I__11074 (
            .O(N__47653),
            .I(N__47473));
    InMux I__11073 (
            .O(N__47650),
            .I(N__47460));
    InMux I__11072 (
            .O(N__47649),
            .I(N__47460));
    InMux I__11071 (
            .O(N__47646),
            .I(N__47460));
    InMux I__11070 (
            .O(N__47645),
            .I(N__47460));
    InMux I__11069 (
            .O(N__47642),
            .I(N__47460));
    InMux I__11068 (
            .O(N__47641),
            .I(N__47460));
    Span12Mux_v I__11067 (
            .O(N__47638),
            .I(N__47455));
    LocalMux I__11066 (
            .O(N__47631),
            .I(N__47455));
    LocalMux I__11065 (
            .O(N__47624),
            .I(N__47452));
    InMux I__11064 (
            .O(N__47623),
            .I(N__47445));
    InMux I__11063 (
            .O(N__47620),
            .I(N__47445));
    InMux I__11062 (
            .O(N__47619),
            .I(N__47445));
    InMux I__11061 (
            .O(N__47618),
            .I(N__47430));
    InMux I__11060 (
            .O(N__47617),
            .I(N__47430));
    InMux I__11059 (
            .O(N__47616),
            .I(N__47430));
    InMux I__11058 (
            .O(N__47615),
            .I(N__47430));
    InMux I__11057 (
            .O(N__47614),
            .I(N__47430));
    InMux I__11056 (
            .O(N__47613),
            .I(N__47430));
    InMux I__11055 (
            .O(N__47612),
            .I(N__47430));
    CascadeMux I__11054 (
            .O(N__47611),
            .I(N__47423));
    CascadeMux I__11053 (
            .O(N__47610),
            .I(N__47420));
    Span4Mux_v I__11052 (
            .O(N__47607),
            .I(N__47407));
    LocalMux I__11051 (
            .O(N__47604),
            .I(N__47407));
    LocalMux I__11050 (
            .O(N__47597),
            .I(N__47407));
    Span4Mux_h I__11049 (
            .O(N__47594),
            .I(N__47407));
    LocalMux I__11048 (
            .O(N__47591),
            .I(N__47407));
    CascadeMux I__11047 (
            .O(N__47590),
            .I(N__47404));
    CascadeMux I__11046 (
            .O(N__47589),
            .I(N__47400));
    CascadeMux I__11045 (
            .O(N__47588),
            .I(N__47396));
    CascadeMux I__11044 (
            .O(N__47587),
            .I(N__47392));
    CascadeMux I__11043 (
            .O(N__47586),
            .I(N__47388));
    CascadeMux I__11042 (
            .O(N__47585),
            .I(N__47384));
    CascadeMux I__11041 (
            .O(N__47584),
            .I(N__47380));
    Span4Mux_h I__11040 (
            .O(N__47579),
            .I(N__47358));
    LocalMux I__11039 (
            .O(N__47564),
            .I(N__47358));
    LocalMux I__11038 (
            .O(N__47547),
            .I(N__47358));
    Span4Mux_h I__11037 (
            .O(N__47542),
            .I(N__47358));
    LocalMux I__11036 (
            .O(N__47527),
            .I(N__47358));
    Span4Mux_v I__11035 (
            .O(N__47524),
            .I(N__47358));
    LocalMux I__11034 (
            .O(N__47507),
            .I(N__47358));
    LocalMux I__11033 (
            .O(N__47490),
            .I(N__47358));
    LocalMux I__11032 (
            .O(N__47473),
            .I(N__47358));
    LocalMux I__11031 (
            .O(N__47460),
            .I(N__47358));
    Span12Mux_s11_h I__11030 (
            .O(N__47455),
            .I(N__47355));
    Span4Mux_h I__11029 (
            .O(N__47452),
            .I(N__47348));
    LocalMux I__11028 (
            .O(N__47445),
            .I(N__47348));
    LocalMux I__11027 (
            .O(N__47430),
            .I(N__47348));
    InMux I__11026 (
            .O(N__47429),
            .I(N__47335));
    InMux I__11025 (
            .O(N__47428),
            .I(N__47335));
    InMux I__11024 (
            .O(N__47427),
            .I(N__47335));
    InMux I__11023 (
            .O(N__47426),
            .I(N__47335));
    InMux I__11022 (
            .O(N__47423),
            .I(N__47335));
    InMux I__11021 (
            .O(N__47420),
            .I(N__47335));
    InMux I__11020 (
            .O(N__47419),
            .I(N__47330));
    InMux I__11019 (
            .O(N__47418),
            .I(N__47330));
    Span4Mux_v I__11018 (
            .O(N__47407),
            .I(N__47327));
    InMux I__11017 (
            .O(N__47404),
            .I(N__47310));
    InMux I__11016 (
            .O(N__47403),
            .I(N__47310));
    InMux I__11015 (
            .O(N__47400),
            .I(N__47310));
    InMux I__11014 (
            .O(N__47399),
            .I(N__47310));
    InMux I__11013 (
            .O(N__47396),
            .I(N__47310));
    InMux I__11012 (
            .O(N__47395),
            .I(N__47310));
    InMux I__11011 (
            .O(N__47392),
            .I(N__47310));
    InMux I__11010 (
            .O(N__47391),
            .I(N__47310));
    InMux I__11009 (
            .O(N__47388),
            .I(N__47297));
    InMux I__11008 (
            .O(N__47387),
            .I(N__47297));
    InMux I__11007 (
            .O(N__47384),
            .I(N__47297));
    InMux I__11006 (
            .O(N__47383),
            .I(N__47297));
    InMux I__11005 (
            .O(N__47380),
            .I(N__47297));
    InMux I__11004 (
            .O(N__47379),
            .I(N__47297));
    Span4Mux_v I__11003 (
            .O(N__47358),
            .I(N__47294));
    Odrv12 I__11002 (
            .O(N__47355),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__11001 (
            .O(N__47348),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11000 (
            .O(N__47335),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10999 (
            .O(N__47330),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10998 (
            .O(N__47327),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10997 (
            .O(N__47310),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10996 (
            .O(N__47297),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10995 (
            .O(N__47294),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__10994 (
            .O(N__47277),
            .I(N__47274));
    LocalMux I__10993 (
            .O(N__47274),
            .I(N__47269));
    InMux I__10992 (
            .O(N__47273),
            .I(N__47266));
    InMux I__10991 (
            .O(N__47272),
            .I(N__47263));
    Span4Mux_v I__10990 (
            .O(N__47269),
            .I(N__47260));
    LocalMux I__10989 (
            .O(N__47266),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__10988 (
            .O(N__47263),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__10987 (
            .O(N__47260),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__10986 (
            .O(N__47253),
            .I(N__47250));
    LocalMux I__10985 (
            .O(N__47250),
            .I(N__47247));
    Odrv12 I__10984 (
            .O(N__47247),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    InMux I__10983 (
            .O(N__47244),
            .I(N__47240));
    CascadeMux I__10982 (
            .O(N__47243),
            .I(N__47237));
    LocalMux I__10981 (
            .O(N__47240),
            .I(N__47234));
    InMux I__10980 (
            .O(N__47237),
            .I(N__47229));
    Span4Mux_h I__10979 (
            .O(N__47234),
            .I(N__47226));
    InMux I__10978 (
            .O(N__47233),
            .I(N__47221));
    InMux I__10977 (
            .O(N__47232),
            .I(N__47221));
    LocalMux I__10976 (
            .O(N__47229),
            .I(N__47218));
    Odrv4 I__10975 (
            .O(N__47226),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__10974 (
            .O(N__47221),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__10973 (
            .O(N__47218),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__10972 (
            .O(N__47211),
            .I(N__47208));
    LocalMux I__10971 (
            .O(N__47208),
            .I(N__47205));
    Span4Mux_h I__10970 (
            .O(N__47205),
            .I(N__47202));
    Span4Mux_h I__10969 (
            .O(N__47202),
            .I(N__47198));
    InMux I__10968 (
            .O(N__47201),
            .I(N__47195));
    Odrv4 I__10967 (
            .O(N__47198),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__10966 (
            .O(N__47195),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__10965 (
            .O(N__47190),
            .I(N__47184));
    InMux I__10964 (
            .O(N__47189),
            .I(N__47184));
    LocalMux I__10963 (
            .O(N__47184),
            .I(N__47181));
    Odrv12 I__10962 (
            .O(N__47181),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__10961 (
            .O(N__47178),
            .I(N__47175));
    InMux I__10960 (
            .O(N__47175),
            .I(N__47169));
    InMux I__10959 (
            .O(N__47174),
            .I(N__47169));
    LocalMux I__10958 (
            .O(N__47169),
            .I(N__47166));
    Odrv12 I__10957 (
            .O(N__47166),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    CEMux I__10956 (
            .O(N__47163),
            .I(N__47127));
    CEMux I__10955 (
            .O(N__47162),
            .I(N__47127));
    CEMux I__10954 (
            .O(N__47161),
            .I(N__47127));
    CEMux I__10953 (
            .O(N__47160),
            .I(N__47127));
    CEMux I__10952 (
            .O(N__47159),
            .I(N__47127));
    CEMux I__10951 (
            .O(N__47158),
            .I(N__47127));
    CEMux I__10950 (
            .O(N__47157),
            .I(N__47127));
    CEMux I__10949 (
            .O(N__47156),
            .I(N__47127));
    CEMux I__10948 (
            .O(N__47155),
            .I(N__47127));
    CEMux I__10947 (
            .O(N__47154),
            .I(N__47127));
    CEMux I__10946 (
            .O(N__47153),
            .I(N__47127));
    CEMux I__10945 (
            .O(N__47152),
            .I(N__47127));
    GlobalMux I__10944 (
            .O(N__47127),
            .I(N__47124));
    gio2CtrlBuf I__10943 (
            .O(N__47124),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    InMux I__10942 (
            .O(N__47121),
            .I(N__47117));
    InMux I__10941 (
            .O(N__47120),
            .I(N__47114));
    LocalMux I__10940 (
            .O(N__47117),
            .I(N__47109));
    LocalMux I__10939 (
            .O(N__47114),
            .I(N__47106));
    InMux I__10938 (
            .O(N__47113),
            .I(N__47103));
    InMux I__10937 (
            .O(N__47112),
            .I(N__47100));
    Span4Mux_v I__10936 (
            .O(N__47109),
            .I(N__47097));
    Span4Mux_v I__10935 (
            .O(N__47106),
            .I(N__47092));
    LocalMux I__10934 (
            .O(N__47103),
            .I(N__47092));
    LocalMux I__10933 (
            .O(N__47100),
            .I(N__47089));
    Span4Mux_h I__10932 (
            .O(N__47097),
            .I(N__47084));
    Span4Mux_h I__10931 (
            .O(N__47092),
            .I(N__47084));
    Span4Mux_v I__10930 (
            .O(N__47089),
            .I(N__47081));
    Odrv4 I__10929 (
            .O(N__47084),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__10928 (
            .O(N__47081),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__10927 (
            .O(N__47076),
            .I(N__47071));
    InMux I__10926 (
            .O(N__47075),
            .I(N__47064));
    InMux I__10925 (
            .O(N__47074),
            .I(N__47064));
    LocalMux I__10924 (
            .O(N__47071),
            .I(N__47061));
    InMux I__10923 (
            .O(N__47070),
            .I(N__47052));
    InMux I__10922 (
            .O(N__47069),
            .I(N__47049));
    LocalMux I__10921 (
            .O(N__47064),
            .I(N__47017));
    Span4Mux_h I__10920 (
            .O(N__47061),
            .I(N__47014));
    InMux I__10919 (
            .O(N__47060),
            .I(N__47007));
    InMux I__10918 (
            .O(N__47059),
            .I(N__47007));
    InMux I__10917 (
            .O(N__47058),
            .I(N__47007));
    InMux I__10916 (
            .O(N__47057),
            .I(N__47000));
    InMux I__10915 (
            .O(N__47056),
            .I(N__47000));
    InMux I__10914 (
            .O(N__47055),
            .I(N__47000));
    LocalMux I__10913 (
            .O(N__47052),
            .I(N__46995));
    LocalMux I__10912 (
            .O(N__47049),
            .I(N__46995));
    InMux I__10911 (
            .O(N__47048),
            .I(N__46992));
    InMux I__10910 (
            .O(N__47047),
            .I(N__46988));
    InMux I__10909 (
            .O(N__47046),
            .I(N__46979));
    InMux I__10908 (
            .O(N__47045),
            .I(N__46979));
    InMux I__10907 (
            .O(N__47044),
            .I(N__46979));
    InMux I__10906 (
            .O(N__47043),
            .I(N__46979));
    InMux I__10905 (
            .O(N__47042),
            .I(N__46972));
    InMux I__10904 (
            .O(N__47041),
            .I(N__46972));
    InMux I__10903 (
            .O(N__47040),
            .I(N__46972));
    CascadeMux I__10902 (
            .O(N__47039),
            .I(N__46966));
    InMux I__10901 (
            .O(N__47038),
            .I(N__46961));
    InMux I__10900 (
            .O(N__47037),
            .I(N__46944));
    InMux I__10899 (
            .O(N__47036),
            .I(N__46944));
    InMux I__10898 (
            .O(N__47035),
            .I(N__46944));
    InMux I__10897 (
            .O(N__47034),
            .I(N__46944));
    InMux I__10896 (
            .O(N__47033),
            .I(N__46944));
    InMux I__10895 (
            .O(N__47032),
            .I(N__46937));
    InMux I__10894 (
            .O(N__47031),
            .I(N__46922));
    InMux I__10893 (
            .O(N__47030),
            .I(N__46922));
    InMux I__10892 (
            .O(N__47029),
            .I(N__46922));
    InMux I__10891 (
            .O(N__47028),
            .I(N__46922));
    InMux I__10890 (
            .O(N__47027),
            .I(N__46922));
    InMux I__10889 (
            .O(N__47026),
            .I(N__46903));
    InMux I__10888 (
            .O(N__47025),
            .I(N__46903));
    InMux I__10887 (
            .O(N__47024),
            .I(N__46903));
    InMux I__10886 (
            .O(N__47023),
            .I(N__46903));
    InMux I__10885 (
            .O(N__47022),
            .I(N__46896));
    InMux I__10884 (
            .O(N__47021),
            .I(N__46896));
    InMux I__10883 (
            .O(N__47020),
            .I(N__46896));
    Span4Mux_h I__10882 (
            .O(N__47017),
            .I(N__46889));
    Span4Mux_v I__10881 (
            .O(N__47014),
            .I(N__46889));
    LocalMux I__10880 (
            .O(N__47007),
            .I(N__46889));
    LocalMux I__10879 (
            .O(N__47000),
            .I(N__46882));
    Span4Mux_v I__10878 (
            .O(N__46995),
            .I(N__46882));
    LocalMux I__10877 (
            .O(N__46992),
            .I(N__46882));
    CascadeMux I__10876 (
            .O(N__46991),
            .I(N__46876));
    LocalMux I__10875 (
            .O(N__46988),
            .I(N__46867));
    LocalMux I__10874 (
            .O(N__46979),
            .I(N__46867));
    LocalMux I__10873 (
            .O(N__46972),
            .I(N__46867));
    InMux I__10872 (
            .O(N__46971),
            .I(N__46854));
    InMux I__10871 (
            .O(N__46970),
            .I(N__46854));
    InMux I__10870 (
            .O(N__46969),
            .I(N__46854));
    InMux I__10869 (
            .O(N__46966),
            .I(N__46854));
    InMux I__10868 (
            .O(N__46965),
            .I(N__46854));
    InMux I__10867 (
            .O(N__46964),
            .I(N__46854));
    LocalMux I__10866 (
            .O(N__46961),
            .I(N__46846));
    InMux I__10865 (
            .O(N__46960),
            .I(N__46835));
    InMux I__10864 (
            .O(N__46959),
            .I(N__46835));
    InMux I__10863 (
            .O(N__46958),
            .I(N__46835));
    InMux I__10862 (
            .O(N__46957),
            .I(N__46835));
    InMux I__10861 (
            .O(N__46956),
            .I(N__46835));
    InMux I__10860 (
            .O(N__46955),
            .I(N__46832));
    LocalMux I__10859 (
            .O(N__46944),
            .I(N__46827));
    InMux I__10858 (
            .O(N__46943),
            .I(N__46818));
    InMux I__10857 (
            .O(N__46942),
            .I(N__46818));
    InMux I__10856 (
            .O(N__46941),
            .I(N__46818));
    InMux I__10855 (
            .O(N__46940),
            .I(N__46818));
    LocalMux I__10854 (
            .O(N__46937),
            .I(N__46808));
    InMux I__10853 (
            .O(N__46936),
            .I(N__46805));
    InMux I__10852 (
            .O(N__46935),
            .I(N__46798));
    InMux I__10851 (
            .O(N__46934),
            .I(N__46798));
    InMux I__10850 (
            .O(N__46933),
            .I(N__46798));
    LocalMux I__10849 (
            .O(N__46922),
            .I(N__46795));
    InMux I__10848 (
            .O(N__46921),
            .I(N__46782));
    InMux I__10847 (
            .O(N__46920),
            .I(N__46782));
    InMux I__10846 (
            .O(N__46919),
            .I(N__46782));
    InMux I__10845 (
            .O(N__46918),
            .I(N__46782));
    InMux I__10844 (
            .O(N__46917),
            .I(N__46782));
    InMux I__10843 (
            .O(N__46916),
            .I(N__46782));
    InMux I__10842 (
            .O(N__46915),
            .I(N__46775));
    InMux I__10841 (
            .O(N__46914),
            .I(N__46775));
    InMux I__10840 (
            .O(N__46913),
            .I(N__46775));
    InMux I__10839 (
            .O(N__46912),
            .I(N__46772));
    LocalMux I__10838 (
            .O(N__46903),
            .I(N__46763));
    LocalMux I__10837 (
            .O(N__46896),
            .I(N__46763));
    Span4Mux_h I__10836 (
            .O(N__46889),
            .I(N__46763));
    Span4Mux_h I__10835 (
            .O(N__46882),
            .I(N__46763));
    InMux I__10834 (
            .O(N__46881),
            .I(N__46760));
    InMux I__10833 (
            .O(N__46880),
            .I(N__46749));
    InMux I__10832 (
            .O(N__46879),
            .I(N__46749));
    InMux I__10831 (
            .O(N__46876),
            .I(N__46749));
    InMux I__10830 (
            .O(N__46875),
            .I(N__46749));
    InMux I__10829 (
            .O(N__46874),
            .I(N__46749));
    Span4Mux_v I__10828 (
            .O(N__46867),
            .I(N__46744));
    LocalMux I__10827 (
            .O(N__46854),
            .I(N__46744));
    InMux I__10826 (
            .O(N__46853),
            .I(N__46733));
    InMux I__10825 (
            .O(N__46852),
            .I(N__46733));
    InMux I__10824 (
            .O(N__46851),
            .I(N__46733));
    InMux I__10823 (
            .O(N__46850),
            .I(N__46733));
    InMux I__10822 (
            .O(N__46849),
            .I(N__46733));
    Span4Mux_h I__10821 (
            .O(N__46846),
            .I(N__46728));
    LocalMux I__10820 (
            .O(N__46835),
            .I(N__46728));
    LocalMux I__10819 (
            .O(N__46832),
            .I(N__46725));
    InMux I__10818 (
            .O(N__46831),
            .I(N__46717));
    InMux I__10817 (
            .O(N__46830),
            .I(N__46717));
    Span4Mux_v I__10816 (
            .O(N__46827),
            .I(N__46712));
    LocalMux I__10815 (
            .O(N__46818),
            .I(N__46712));
    InMux I__10814 (
            .O(N__46817),
            .I(N__46703));
    InMux I__10813 (
            .O(N__46816),
            .I(N__46703));
    InMux I__10812 (
            .O(N__46815),
            .I(N__46703));
    InMux I__10811 (
            .O(N__46814),
            .I(N__46703));
    InMux I__10810 (
            .O(N__46813),
            .I(N__46696));
    InMux I__10809 (
            .O(N__46812),
            .I(N__46696));
    InMux I__10808 (
            .O(N__46811),
            .I(N__46696));
    Span4Mux_v I__10807 (
            .O(N__46808),
            .I(N__46689));
    LocalMux I__10806 (
            .O(N__46805),
            .I(N__46689));
    LocalMux I__10805 (
            .O(N__46798),
            .I(N__46689));
    Span4Mux_h I__10804 (
            .O(N__46795),
            .I(N__46686));
    LocalMux I__10803 (
            .O(N__46782),
            .I(N__46681));
    LocalMux I__10802 (
            .O(N__46775),
            .I(N__46681));
    LocalMux I__10801 (
            .O(N__46772),
            .I(N__46676));
    Span4Mux_v I__10800 (
            .O(N__46763),
            .I(N__46676));
    LocalMux I__10799 (
            .O(N__46760),
            .I(N__46671));
    LocalMux I__10798 (
            .O(N__46749),
            .I(N__46671));
    Span4Mux_h I__10797 (
            .O(N__46744),
            .I(N__46664));
    LocalMux I__10796 (
            .O(N__46733),
            .I(N__46664));
    Span4Mux_v I__10795 (
            .O(N__46728),
            .I(N__46664));
    Span4Mux_h I__10794 (
            .O(N__46725),
            .I(N__46661));
    InMux I__10793 (
            .O(N__46724),
            .I(N__46658));
    InMux I__10792 (
            .O(N__46723),
            .I(N__46653));
    InMux I__10791 (
            .O(N__46722),
            .I(N__46653));
    LocalMux I__10790 (
            .O(N__46717),
            .I(N__46648));
    Span4Mux_v I__10789 (
            .O(N__46712),
            .I(N__46648));
    LocalMux I__10788 (
            .O(N__46703),
            .I(N__46639));
    LocalMux I__10787 (
            .O(N__46696),
            .I(N__46639));
    Span4Mux_h I__10786 (
            .O(N__46689),
            .I(N__46639));
    Span4Mux_v I__10785 (
            .O(N__46686),
            .I(N__46639));
    Span4Mux_v I__10784 (
            .O(N__46681),
            .I(N__46634));
    Span4Mux_h I__10783 (
            .O(N__46676),
            .I(N__46634));
    Span4Mux_h I__10782 (
            .O(N__46671),
            .I(N__46629));
    Span4Mux_v I__10781 (
            .O(N__46664),
            .I(N__46629));
    Span4Mux_v I__10780 (
            .O(N__46661),
            .I(N__46626));
    LocalMux I__10779 (
            .O(N__46658),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__10778 (
            .O(N__46653),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__10777 (
            .O(N__46648),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__10776 (
            .O(N__46639),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__10775 (
            .O(N__46634),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__10774 (
            .O(N__46629),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__10773 (
            .O(N__46626),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__10772 (
            .O(N__46611),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__10771 (
            .O(N__46608),
            .I(N__46605));
    LocalMux I__10770 (
            .O(N__46605),
            .I(N__46601));
    InMux I__10769 (
            .O(N__46604),
            .I(N__46598));
    Span4Mux_h I__10768 (
            .O(N__46601),
            .I(N__46595));
    LocalMux I__10767 (
            .O(N__46598),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__10766 (
            .O(N__46595),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    InMux I__10765 (
            .O(N__46590),
            .I(N__46587));
    LocalMux I__10764 (
            .O(N__46587),
            .I(N__46584));
    Span4Mux_h I__10763 (
            .O(N__46584),
            .I(N__46581));
    Odrv4 I__10762 (
            .O(N__46581),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    CascadeMux I__10761 (
            .O(N__46578),
            .I(N__46573));
    InMux I__10760 (
            .O(N__46577),
            .I(N__46570));
    InMux I__10759 (
            .O(N__46576),
            .I(N__46567));
    InMux I__10758 (
            .O(N__46573),
            .I(N__46564));
    LocalMux I__10757 (
            .O(N__46570),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__10756 (
            .O(N__46567),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__10755 (
            .O(N__46564),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    CascadeMux I__10754 (
            .O(N__46557),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    CascadeMux I__10753 (
            .O(N__46554),
            .I(N__46550));
    InMux I__10752 (
            .O(N__46553),
            .I(N__46547));
    InMux I__10751 (
            .O(N__46550),
            .I(N__46544));
    LocalMux I__10750 (
            .O(N__46547),
            .I(N__46539));
    LocalMux I__10749 (
            .O(N__46544),
            .I(N__46539));
    Span4Mux_h I__10748 (
            .O(N__46539),
            .I(N__46536));
    Span4Mux_v I__10747 (
            .O(N__46536),
            .I(N__46533));
    Odrv4 I__10746 (
            .O(N__46533),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__10745 (
            .O(N__46530),
            .I(N__46526));
    InMux I__10744 (
            .O(N__46529),
            .I(N__46522));
    LocalMux I__10743 (
            .O(N__46526),
            .I(N__46519));
    InMux I__10742 (
            .O(N__46525),
            .I(N__46516));
    LocalMux I__10741 (
            .O(N__46522),
            .I(N__46513));
    Span4Mux_v I__10740 (
            .O(N__46519),
            .I(N__46510));
    LocalMux I__10739 (
            .O(N__46516),
            .I(N__46507));
    Span12Mux_v I__10738 (
            .O(N__46513),
            .I(N__46504));
    Span4Mux_v I__10737 (
            .O(N__46510),
            .I(N__46499));
    Span4Mux_v I__10736 (
            .O(N__46507),
            .I(N__46499));
    Odrv12 I__10735 (
            .O(N__46504),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__10734 (
            .O(N__46499),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__10733 (
            .O(N__46494),
            .I(N__46491));
    LocalMux I__10732 (
            .O(N__46491),
            .I(N__46487));
    InMux I__10731 (
            .O(N__46490),
            .I(N__46484));
    Span4Mux_h I__10730 (
            .O(N__46487),
            .I(N__46480));
    LocalMux I__10729 (
            .O(N__46484),
            .I(N__46477));
    InMux I__10728 (
            .O(N__46483),
            .I(N__46474));
    Span4Mux_v I__10727 (
            .O(N__46480),
            .I(N__46469));
    Span4Mux_h I__10726 (
            .O(N__46477),
            .I(N__46469));
    LocalMux I__10725 (
            .O(N__46474),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__10724 (
            .O(N__46469),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__10723 (
            .O(N__46464),
            .I(N__46461));
    LocalMux I__10722 (
            .O(N__46461),
            .I(N__46455));
    InMux I__10721 (
            .O(N__46460),
            .I(N__46452));
    InMux I__10720 (
            .O(N__46459),
            .I(N__46447));
    InMux I__10719 (
            .O(N__46458),
            .I(N__46447));
    Odrv4 I__10718 (
            .O(N__46455),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__10717 (
            .O(N__46452),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__10716 (
            .O(N__46447),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    InMux I__10715 (
            .O(N__46440),
            .I(N__46436));
    InMux I__10714 (
            .O(N__46439),
            .I(N__46433));
    LocalMux I__10713 (
            .O(N__46436),
            .I(N__46429));
    LocalMux I__10712 (
            .O(N__46433),
            .I(N__46426));
    InMux I__10711 (
            .O(N__46432),
            .I(N__46423));
    Span4Mux_v I__10710 (
            .O(N__46429),
            .I(N__46418));
    Span4Mux_h I__10709 (
            .O(N__46426),
            .I(N__46418));
    LocalMux I__10708 (
            .O(N__46423),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__10707 (
            .O(N__46418),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    CEMux I__10706 (
            .O(N__46413),
            .I(N__46389));
    CEMux I__10705 (
            .O(N__46412),
            .I(N__46389));
    CEMux I__10704 (
            .O(N__46411),
            .I(N__46389));
    CEMux I__10703 (
            .O(N__46410),
            .I(N__46389));
    CEMux I__10702 (
            .O(N__46409),
            .I(N__46389));
    CEMux I__10701 (
            .O(N__46408),
            .I(N__46389));
    CEMux I__10700 (
            .O(N__46407),
            .I(N__46389));
    CEMux I__10699 (
            .O(N__46406),
            .I(N__46389));
    GlobalMux I__10698 (
            .O(N__46389),
            .I(N__46386));
    gio2CtrlBuf I__10697 (
            .O(N__46386),
            .I(\current_shift_inst.timer_s1.N_161_i_g ));
    InMux I__10696 (
            .O(N__46383),
            .I(N__46380));
    LocalMux I__10695 (
            .O(N__46380),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__10694 (
            .O(N__46377),
            .I(N__46373));
    CascadeMux I__10693 (
            .O(N__46376),
            .I(N__46370));
    InMux I__10692 (
            .O(N__46373),
            .I(N__46366));
    InMux I__10691 (
            .O(N__46370),
            .I(N__46363));
    InMux I__10690 (
            .O(N__46369),
            .I(N__46360));
    LocalMux I__10689 (
            .O(N__46366),
            .I(N__46354));
    LocalMux I__10688 (
            .O(N__46363),
            .I(N__46354));
    LocalMux I__10687 (
            .O(N__46360),
            .I(N__46351));
    InMux I__10686 (
            .O(N__46359),
            .I(N__46348));
    Span4Mux_v I__10685 (
            .O(N__46354),
            .I(N__46343));
    Span4Mux_v I__10684 (
            .O(N__46351),
            .I(N__46343));
    LocalMux I__10683 (
            .O(N__46348),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__10682 (
            .O(N__46343),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__10681 (
            .O(N__46338),
            .I(N__46335));
    InMux I__10680 (
            .O(N__46335),
            .I(N__46332));
    LocalMux I__10679 (
            .O(N__46332),
            .I(N__46329));
    Odrv12 I__10678 (
            .O(N__46329),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__10677 (
            .O(N__46326),
            .I(N__46323));
    InMux I__10676 (
            .O(N__46323),
            .I(N__46319));
    InMux I__10675 (
            .O(N__46322),
            .I(N__46316));
    LocalMux I__10674 (
            .O(N__46319),
            .I(N__46310));
    LocalMux I__10673 (
            .O(N__46316),
            .I(N__46310));
    InMux I__10672 (
            .O(N__46315),
            .I(N__46307));
    Span4Mux_h I__10671 (
            .O(N__46310),
            .I(N__46304));
    LocalMux I__10670 (
            .O(N__46307),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__10669 (
            .O(N__46304),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__10668 (
            .O(N__46299),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    CascadeMux I__10667 (
            .O(N__46296),
            .I(N__46293));
    InMux I__10666 (
            .O(N__46293),
            .I(N__46289));
    InMux I__10665 (
            .O(N__46292),
            .I(N__46286));
    LocalMux I__10664 (
            .O(N__46289),
            .I(N__46280));
    LocalMux I__10663 (
            .O(N__46286),
            .I(N__46280));
    InMux I__10662 (
            .O(N__46285),
            .I(N__46277));
    Span4Mux_v I__10661 (
            .O(N__46280),
            .I(N__46274));
    LocalMux I__10660 (
            .O(N__46277),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__10659 (
            .O(N__46274),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__10658 (
            .O(N__46269),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__10657 (
            .O(N__46266),
            .I(N__46260));
    InMux I__10656 (
            .O(N__46265),
            .I(N__46260));
    LocalMux I__10655 (
            .O(N__46260),
            .I(N__46256));
    InMux I__10654 (
            .O(N__46259),
            .I(N__46253));
    Span4Mux_h I__10653 (
            .O(N__46256),
            .I(N__46250));
    LocalMux I__10652 (
            .O(N__46253),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__10651 (
            .O(N__46250),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__10650 (
            .O(N__46245),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__10649 (
            .O(N__46242),
            .I(N__46239));
    InMux I__10648 (
            .O(N__46239),
            .I(N__46234));
    InMux I__10647 (
            .O(N__46238),
            .I(N__46231));
    InMux I__10646 (
            .O(N__46237),
            .I(N__46228));
    LocalMux I__10645 (
            .O(N__46234),
            .I(N__46225));
    LocalMux I__10644 (
            .O(N__46231),
            .I(N__46222));
    LocalMux I__10643 (
            .O(N__46228),
            .I(N__46217));
    Span4Mux_v I__10642 (
            .O(N__46225),
            .I(N__46217));
    Span4Mux_h I__10641 (
            .O(N__46222),
            .I(N__46214));
    Odrv4 I__10640 (
            .O(N__46217),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__10639 (
            .O(N__46214),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__10638 (
            .O(N__46209),
            .I(bfn_18_14_0_));
    CascadeMux I__10637 (
            .O(N__46206),
            .I(N__46202));
    CascadeMux I__10636 (
            .O(N__46205),
            .I(N__46199));
    InMux I__10635 (
            .O(N__46202),
            .I(N__46196));
    InMux I__10634 (
            .O(N__46199),
            .I(N__46193));
    LocalMux I__10633 (
            .O(N__46196),
            .I(N__46189));
    LocalMux I__10632 (
            .O(N__46193),
            .I(N__46186));
    InMux I__10631 (
            .O(N__46192),
            .I(N__46183));
    Span4Mux_v I__10630 (
            .O(N__46189),
            .I(N__46180));
    Span4Mux_h I__10629 (
            .O(N__46186),
            .I(N__46177));
    LocalMux I__10628 (
            .O(N__46183),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__10627 (
            .O(N__46180),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__10626 (
            .O(N__46177),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__10625 (
            .O(N__46170),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__10624 (
            .O(N__46167),
            .I(N__46161));
    InMux I__10623 (
            .O(N__46166),
            .I(N__46161));
    LocalMux I__10622 (
            .O(N__46161),
            .I(N__46157));
    InMux I__10621 (
            .O(N__46160),
            .I(N__46154));
    Span4Mux_h I__10620 (
            .O(N__46157),
            .I(N__46151));
    LocalMux I__10619 (
            .O(N__46154),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv4 I__10618 (
            .O(N__46151),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__10617 (
            .O(N__46146),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__10616 (
            .O(N__46143),
            .I(N__46140));
    InMux I__10615 (
            .O(N__46140),
            .I(N__46136));
    InMux I__10614 (
            .O(N__46139),
            .I(N__46133));
    LocalMux I__10613 (
            .O(N__46136),
            .I(N__46127));
    LocalMux I__10612 (
            .O(N__46133),
            .I(N__46127));
    InMux I__10611 (
            .O(N__46132),
            .I(N__46124));
    Span4Mux_h I__10610 (
            .O(N__46127),
            .I(N__46121));
    LocalMux I__10609 (
            .O(N__46124),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv4 I__10608 (
            .O(N__46121),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__10607 (
            .O(N__46116),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    CascadeMux I__10606 (
            .O(N__46113),
            .I(N__46110));
    InMux I__10605 (
            .O(N__46110),
            .I(N__46107));
    LocalMux I__10604 (
            .O(N__46107),
            .I(N__46103));
    InMux I__10603 (
            .O(N__46106),
            .I(N__46100));
    Span4Mux_h I__10602 (
            .O(N__46103),
            .I(N__46097));
    LocalMux I__10601 (
            .O(N__46100),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__10600 (
            .O(N__46097),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__10599 (
            .O(N__46092),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    CascadeMux I__10598 (
            .O(N__46089),
            .I(N__46086));
    InMux I__10597 (
            .O(N__46086),
            .I(N__46082));
    InMux I__10596 (
            .O(N__46085),
            .I(N__46079));
    LocalMux I__10595 (
            .O(N__46082),
            .I(N__46073));
    LocalMux I__10594 (
            .O(N__46079),
            .I(N__46073));
    InMux I__10593 (
            .O(N__46078),
            .I(N__46070));
    Span4Mux_h I__10592 (
            .O(N__46073),
            .I(N__46067));
    LocalMux I__10591 (
            .O(N__46070),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__10590 (
            .O(N__46067),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__10589 (
            .O(N__46062),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__10588 (
            .O(N__46059),
            .I(N__46055));
    CascadeMux I__10587 (
            .O(N__46058),
            .I(N__46052));
    InMux I__10586 (
            .O(N__46055),
            .I(N__46047));
    InMux I__10585 (
            .O(N__46052),
            .I(N__46047));
    LocalMux I__10584 (
            .O(N__46047),
            .I(N__46043));
    InMux I__10583 (
            .O(N__46046),
            .I(N__46040));
    Span4Mux_h I__10582 (
            .O(N__46043),
            .I(N__46037));
    LocalMux I__10581 (
            .O(N__46040),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__10580 (
            .O(N__46037),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__10579 (
            .O(N__46032),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    CascadeMux I__10578 (
            .O(N__46029),
            .I(N__46026));
    InMux I__10577 (
            .O(N__46026),
            .I(N__46022));
    InMux I__10576 (
            .O(N__46025),
            .I(N__46019));
    LocalMux I__10575 (
            .O(N__46022),
            .I(N__46013));
    LocalMux I__10574 (
            .O(N__46019),
            .I(N__46013));
    InMux I__10573 (
            .O(N__46018),
            .I(N__46010));
    Span4Mux_h I__10572 (
            .O(N__46013),
            .I(N__46007));
    LocalMux I__10571 (
            .O(N__46010),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__10570 (
            .O(N__46007),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__10569 (
            .O(N__46002),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__10568 (
            .O(N__45999),
            .I(N__45992));
    InMux I__10567 (
            .O(N__45998),
            .I(N__45992));
    InMux I__10566 (
            .O(N__45997),
            .I(N__45989));
    LocalMux I__10565 (
            .O(N__45992),
            .I(N__45986));
    LocalMux I__10564 (
            .O(N__45989),
            .I(N__45981));
    Span4Mux_v I__10563 (
            .O(N__45986),
            .I(N__45981));
    Odrv4 I__10562 (
            .O(N__45981),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__10561 (
            .O(N__45978),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__10560 (
            .O(N__45975),
            .I(N__45972));
    InMux I__10559 (
            .O(N__45972),
            .I(N__45968));
    InMux I__10558 (
            .O(N__45971),
            .I(N__45965));
    LocalMux I__10557 (
            .O(N__45968),
            .I(N__45961));
    LocalMux I__10556 (
            .O(N__45965),
            .I(N__45958));
    InMux I__10555 (
            .O(N__45964),
            .I(N__45955));
    Span4Mux_v I__10554 (
            .O(N__45961),
            .I(N__45952));
    Span4Mux_h I__10553 (
            .O(N__45958),
            .I(N__45949));
    LocalMux I__10552 (
            .O(N__45955),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__10551 (
            .O(N__45952),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__10550 (
            .O(N__45949),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__10549 (
            .O(N__45942),
            .I(bfn_18_13_0_));
    CascadeMux I__10548 (
            .O(N__45939),
            .I(N__45935));
    CascadeMux I__10547 (
            .O(N__45938),
            .I(N__45932));
    InMux I__10546 (
            .O(N__45935),
            .I(N__45929));
    InMux I__10545 (
            .O(N__45932),
            .I(N__45926));
    LocalMux I__10544 (
            .O(N__45929),
            .I(N__45920));
    LocalMux I__10543 (
            .O(N__45926),
            .I(N__45920));
    InMux I__10542 (
            .O(N__45925),
            .I(N__45917));
    Span4Mux_v I__10541 (
            .O(N__45920),
            .I(N__45914));
    LocalMux I__10540 (
            .O(N__45917),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__10539 (
            .O(N__45914),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__10538 (
            .O(N__45909),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__10537 (
            .O(N__45906),
            .I(N__45903));
    InMux I__10536 (
            .O(N__45903),
            .I(N__45899));
    InMux I__10535 (
            .O(N__45902),
            .I(N__45896));
    LocalMux I__10534 (
            .O(N__45899),
            .I(N__45890));
    LocalMux I__10533 (
            .O(N__45896),
            .I(N__45890));
    InMux I__10532 (
            .O(N__45895),
            .I(N__45887));
    Span4Mux_h I__10531 (
            .O(N__45890),
            .I(N__45884));
    LocalMux I__10530 (
            .O(N__45887),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__10529 (
            .O(N__45884),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__10528 (
            .O(N__45879),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__10527 (
            .O(N__45876),
            .I(N__45873));
    InMux I__10526 (
            .O(N__45873),
            .I(N__45869));
    InMux I__10525 (
            .O(N__45872),
            .I(N__45866));
    LocalMux I__10524 (
            .O(N__45869),
            .I(N__45860));
    LocalMux I__10523 (
            .O(N__45866),
            .I(N__45860));
    InMux I__10522 (
            .O(N__45865),
            .I(N__45857));
    Span4Mux_h I__10521 (
            .O(N__45860),
            .I(N__45854));
    LocalMux I__10520 (
            .O(N__45857),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv4 I__10519 (
            .O(N__45854),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__10518 (
            .O(N__45849),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    CascadeMux I__10517 (
            .O(N__45846),
            .I(N__45843));
    InMux I__10516 (
            .O(N__45843),
            .I(N__45839));
    InMux I__10515 (
            .O(N__45842),
            .I(N__45836));
    LocalMux I__10514 (
            .O(N__45839),
            .I(N__45830));
    LocalMux I__10513 (
            .O(N__45836),
            .I(N__45830));
    InMux I__10512 (
            .O(N__45835),
            .I(N__45827));
    Span4Mux_h I__10511 (
            .O(N__45830),
            .I(N__45824));
    LocalMux I__10510 (
            .O(N__45827),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__10509 (
            .O(N__45824),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__10508 (
            .O(N__45819),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__10507 (
            .O(N__45816),
            .I(N__45812));
    CascadeMux I__10506 (
            .O(N__45815),
            .I(N__45809));
    InMux I__10505 (
            .O(N__45812),
            .I(N__45804));
    InMux I__10504 (
            .O(N__45809),
            .I(N__45804));
    LocalMux I__10503 (
            .O(N__45804),
            .I(N__45800));
    InMux I__10502 (
            .O(N__45803),
            .I(N__45797));
    Span4Mux_h I__10501 (
            .O(N__45800),
            .I(N__45794));
    LocalMux I__10500 (
            .O(N__45797),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__10499 (
            .O(N__45794),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__10498 (
            .O(N__45789),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__10497 (
            .O(N__45786),
            .I(N__45782));
    CascadeMux I__10496 (
            .O(N__45785),
            .I(N__45779));
    InMux I__10495 (
            .O(N__45782),
            .I(N__45774));
    InMux I__10494 (
            .O(N__45779),
            .I(N__45774));
    LocalMux I__10493 (
            .O(N__45774),
            .I(N__45770));
    InMux I__10492 (
            .O(N__45773),
            .I(N__45767));
    Span4Mux_h I__10491 (
            .O(N__45770),
            .I(N__45764));
    LocalMux I__10490 (
            .O(N__45767),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__10489 (
            .O(N__45764),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__10488 (
            .O(N__45759),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__10487 (
            .O(N__45756),
            .I(N__45750));
    InMux I__10486 (
            .O(N__45755),
            .I(N__45750));
    LocalMux I__10485 (
            .O(N__45750),
            .I(N__45746));
    InMux I__10484 (
            .O(N__45749),
            .I(N__45743));
    Span4Mux_h I__10483 (
            .O(N__45746),
            .I(N__45740));
    LocalMux I__10482 (
            .O(N__45743),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__10481 (
            .O(N__45740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__10480 (
            .O(N__45735),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__10479 (
            .O(N__45732),
            .I(N__45726));
    InMux I__10478 (
            .O(N__45731),
            .I(N__45726));
    LocalMux I__10477 (
            .O(N__45726),
            .I(N__45722));
    InMux I__10476 (
            .O(N__45725),
            .I(N__45719));
    Span4Mux_h I__10475 (
            .O(N__45722),
            .I(N__45716));
    LocalMux I__10474 (
            .O(N__45719),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__10473 (
            .O(N__45716),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__10472 (
            .O(N__45711),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__10471 (
            .O(N__45708),
            .I(N__45704));
    CascadeMux I__10470 (
            .O(N__45707),
            .I(N__45701));
    InMux I__10469 (
            .O(N__45704),
            .I(N__45698));
    InMux I__10468 (
            .O(N__45701),
            .I(N__45695));
    LocalMux I__10467 (
            .O(N__45698),
            .I(N__45691));
    LocalMux I__10466 (
            .O(N__45695),
            .I(N__45688));
    InMux I__10465 (
            .O(N__45694),
            .I(N__45685));
    Span4Mux_v I__10464 (
            .O(N__45691),
            .I(N__45682));
    Span4Mux_h I__10463 (
            .O(N__45688),
            .I(N__45679));
    LocalMux I__10462 (
            .O(N__45685),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__10461 (
            .O(N__45682),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__10460 (
            .O(N__45679),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__10459 (
            .O(N__45672),
            .I(bfn_18_12_0_));
    CascadeMux I__10458 (
            .O(N__45669),
            .I(N__45665));
    CascadeMux I__10457 (
            .O(N__45668),
            .I(N__45662));
    InMux I__10456 (
            .O(N__45665),
            .I(N__45659));
    InMux I__10455 (
            .O(N__45662),
            .I(N__45656));
    LocalMux I__10454 (
            .O(N__45659),
            .I(N__45652));
    LocalMux I__10453 (
            .O(N__45656),
            .I(N__45649));
    InMux I__10452 (
            .O(N__45655),
            .I(N__45646));
    Span4Mux_v I__10451 (
            .O(N__45652),
            .I(N__45643));
    Span4Mux_h I__10450 (
            .O(N__45649),
            .I(N__45640));
    LocalMux I__10449 (
            .O(N__45646),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__10448 (
            .O(N__45643),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__10447 (
            .O(N__45640),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__10446 (
            .O(N__45633),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__10445 (
            .O(N__45630),
            .I(N__45627));
    InMux I__10444 (
            .O(N__45627),
            .I(N__45623));
    InMux I__10443 (
            .O(N__45626),
            .I(N__45620));
    LocalMux I__10442 (
            .O(N__45623),
            .I(N__45614));
    LocalMux I__10441 (
            .O(N__45620),
            .I(N__45614));
    InMux I__10440 (
            .O(N__45619),
            .I(N__45611));
    Span4Mux_h I__10439 (
            .O(N__45614),
            .I(N__45608));
    LocalMux I__10438 (
            .O(N__45611),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__10437 (
            .O(N__45608),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__10436 (
            .O(N__45603),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__10435 (
            .O(N__45600),
            .I(N__45594));
    InMux I__10434 (
            .O(N__45599),
            .I(N__45594));
    LocalMux I__10433 (
            .O(N__45594),
            .I(N__45590));
    InMux I__10432 (
            .O(N__45593),
            .I(N__45587));
    Span4Mux_h I__10431 (
            .O(N__45590),
            .I(N__45584));
    LocalMux I__10430 (
            .O(N__45587),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__10429 (
            .O(N__45584),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__10428 (
            .O(N__45579),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__10427 (
            .O(N__45576),
            .I(N__45570));
    InMux I__10426 (
            .O(N__45575),
            .I(N__45570));
    LocalMux I__10425 (
            .O(N__45570),
            .I(N__45567));
    Odrv12 I__10424 (
            .O(N__45567),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    CascadeMux I__10423 (
            .O(N__45564),
            .I(N__45559));
    InMux I__10422 (
            .O(N__45563),
            .I(N__45556));
    InMux I__10421 (
            .O(N__45562),
            .I(N__45551));
    InMux I__10420 (
            .O(N__45559),
            .I(N__45551));
    LocalMux I__10419 (
            .O(N__45556),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__10418 (
            .O(N__45551),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__10417 (
            .O(N__45546),
            .I(N__45541));
    InMux I__10416 (
            .O(N__45545),
            .I(N__45536));
    InMux I__10415 (
            .O(N__45544),
            .I(N__45536));
    LocalMux I__10414 (
            .O(N__45541),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    LocalMux I__10413 (
            .O(N__45536),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    CascadeMux I__10412 (
            .O(N__45531),
            .I(N__45528));
    InMux I__10411 (
            .O(N__45528),
            .I(N__45525));
    LocalMux I__10410 (
            .O(N__45525),
            .I(N__45522));
    Span4Mux_v I__10409 (
            .O(N__45522),
            .I(N__45519));
    Odrv4 I__10408 (
            .O(N__45519),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    CascadeMux I__10407 (
            .O(N__45516),
            .I(N__45511));
    InMux I__10406 (
            .O(N__45515),
            .I(N__45508));
    CascadeMux I__10405 (
            .O(N__45514),
            .I(N__45504));
    InMux I__10404 (
            .O(N__45511),
            .I(N__45501));
    LocalMux I__10403 (
            .O(N__45508),
            .I(N__45498));
    InMux I__10402 (
            .O(N__45507),
            .I(N__45493));
    InMux I__10401 (
            .O(N__45504),
            .I(N__45493));
    LocalMux I__10400 (
            .O(N__45501),
            .I(N__45490));
    Span4Mux_v I__10399 (
            .O(N__45498),
            .I(N__45487));
    LocalMux I__10398 (
            .O(N__45493),
            .I(N__45484));
    Span4Mux_h I__10397 (
            .O(N__45490),
            .I(N__45481));
    Odrv4 I__10396 (
            .O(N__45487),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__10395 (
            .O(N__45484),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__10394 (
            .O(N__45481),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__10393 (
            .O(N__45474),
            .I(N__45471));
    LocalMux I__10392 (
            .O(N__45471),
            .I(N__45468));
    Span4Mux_h I__10391 (
            .O(N__45468),
            .I(N__45464));
    InMux I__10390 (
            .O(N__45467),
            .I(N__45461));
    Odrv4 I__10389 (
            .O(N__45464),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    LocalMux I__10388 (
            .O(N__45461),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    CascadeMux I__10387 (
            .O(N__45456),
            .I(N__45452));
    InMux I__10386 (
            .O(N__45455),
            .I(N__45447));
    InMux I__10385 (
            .O(N__45452),
            .I(N__45447));
    LocalMux I__10384 (
            .O(N__45447),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    InMux I__10383 (
            .O(N__45444),
            .I(N__45436));
    InMux I__10382 (
            .O(N__45443),
            .I(N__45436));
    InMux I__10381 (
            .O(N__45442),
            .I(N__45433));
    InMux I__10380 (
            .O(N__45441),
            .I(N__45430));
    LocalMux I__10379 (
            .O(N__45436),
            .I(N__45425));
    LocalMux I__10378 (
            .O(N__45433),
            .I(N__45425));
    LocalMux I__10377 (
            .O(N__45430),
            .I(N__45422));
    Span4Mux_v I__10376 (
            .O(N__45425),
            .I(N__45419));
    Odrv12 I__10375 (
            .O(N__45422),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv4 I__10374 (
            .O(N__45419),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__10373 (
            .O(N__45414),
            .I(N__45411));
    LocalMux I__10372 (
            .O(N__45411),
            .I(N__45408));
    Span12Mux_s10_v I__10371 (
            .O(N__45408),
            .I(N__45404));
    InMux I__10370 (
            .O(N__45407),
            .I(N__45401));
    Odrv12 I__10369 (
            .O(N__45404),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    LocalMux I__10368 (
            .O(N__45401),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    InMux I__10367 (
            .O(N__45396),
            .I(N__45393));
    LocalMux I__10366 (
            .O(N__45393),
            .I(N__45390));
    Span4Mux_v I__10365 (
            .O(N__45390),
            .I(N__45387));
    Odrv4 I__10364 (
            .O(N__45387),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    InMux I__10363 (
            .O(N__45384),
            .I(N__45380));
    InMux I__10362 (
            .O(N__45383),
            .I(N__45377));
    LocalMux I__10361 (
            .O(N__45380),
            .I(N__45373));
    LocalMux I__10360 (
            .O(N__45377),
            .I(N__45370));
    InMux I__10359 (
            .O(N__45376),
            .I(N__45367));
    Span4Mux_h I__10358 (
            .O(N__45373),
            .I(N__45364));
    Span4Mux_h I__10357 (
            .O(N__45370),
            .I(N__45361));
    LocalMux I__10356 (
            .O(N__45367),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    Odrv4 I__10355 (
            .O(N__45364),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    Odrv4 I__10354 (
            .O(N__45361),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    InMux I__10353 (
            .O(N__45354),
            .I(N__45349));
    InMux I__10352 (
            .O(N__45353),
            .I(N__45346));
    InMux I__10351 (
            .O(N__45352),
            .I(N__45343));
    LocalMux I__10350 (
            .O(N__45349),
            .I(N__45337));
    LocalMux I__10349 (
            .O(N__45346),
            .I(N__45337));
    LocalMux I__10348 (
            .O(N__45343),
            .I(N__45334));
    InMux I__10347 (
            .O(N__45342),
            .I(N__45331));
    Span4Mux_v I__10346 (
            .O(N__45337),
            .I(N__45328));
    Odrv4 I__10345 (
            .O(N__45334),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    LocalMux I__10344 (
            .O(N__45331),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__10343 (
            .O(N__45328),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__10342 (
            .O(N__45321),
            .I(N__45318));
    LocalMux I__10341 (
            .O(N__45318),
            .I(N__45315));
    Span4Mux_v I__10340 (
            .O(N__45315),
            .I(N__45312));
    Odrv4 I__10339 (
            .O(N__45312),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__10338 (
            .O(N__45309),
            .I(bfn_18_11_0_));
    CascadeMux I__10337 (
            .O(N__45306),
            .I(N__45302));
    InMux I__10336 (
            .O(N__45305),
            .I(N__45299));
    InMux I__10335 (
            .O(N__45302),
            .I(N__45296));
    LocalMux I__10334 (
            .O(N__45299),
            .I(N__45292));
    LocalMux I__10333 (
            .O(N__45296),
            .I(N__45289));
    InMux I__10332 (
            .O(N__45295),
            .I(N__45286));
    Span4Mux_v I__10331 (
            .O(N__45292),
            .I(N__45281));
    Span4Mux_v I__10330 (
            .O(N__45289),
            .I(N__45281));
    LocalMux I__10329 (
            .O(N__45286),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__10328 (
            .O(N__45281),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__10327 (
            .O(N__45276),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__10326 (
            .O(N__45273),
            .I(N__45267));
    InMux I__10325 (
            .O(N__45272),
            .I(N__45267));
    LocalMux I__10324 (
            .O(N__45267),
            .I(N__45263));
    InMux I__10323 (
            .O(N__45266),
            .I(N__45260));
    Span4Mux_h I__10322 (
            .O(N__45263),
            .I(N__45257));
    LocalMux I__10321 (
            .O(N__45260),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__10320 (
            .O(N__45257),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__10319 (
            .O(N__45252),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__10318 (
            .O(N__45249),
            .I(N__45243));
    InMux I__10317 (
            .O(N__45248),
            .I(N__45243));
    LocalMux I__10316 (
            .O(N__45243),
            .I(N__45239));
    InMux I__10315 (
            .O(N__45242),
            .I(N__45236));
    Span4Mux_h I__10314 (
            .O(N__45239),
            .I(N__45233));
    LocalMux I__10313 (
            .O(N__45236),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__10312 (
            .O(N__45233),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__10311 (
            .O(N__45228),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__10310 (
            .O(N__45225),
            .I(N__45222));
    LocalMux I__10309 (
            .O(N__45222),
            .I(N__45219));
    Odrv4 I__10308 (
            .O(N__45219),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__10307 (
            .O(N__45216),
            .I(N__45213));
    LocalMux I__10306 (
            .O(N__45213),
            .I(N__45209));
    InMux I__10305 (
            .O(N__45212),
            .I(N__45205));
    Span4Mux_h I__10304 (
            .O(N__45209),
            .I(N__45202));
    InMux I__10303 (
            .O(N__45208),
            .I(N__45199));
    LocalMux I__10302 (
            .O(N__45205),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    Odrv4 I__10301 (
            .O(N__45202),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__10300 (
            .O(N__45199),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__10299 (
            .O(N__45192),
            .I(N__45187));
    InMux I__10298 (
            .O(N__45191),
            .I(N__45184));
    InMux I__10297 (
            .O(N__45190),
            .I(N__45181));
    LocalMux I__10296 (
            .O(N__45187),
            .I(N__45178));
    LocalMux I__10295 (
            .O(N__45184),
            .I(N__45173));
    LocalMux I__10294 (
            .O(N__45181),
            .I(N__45173));
    Span4Mux_v I__10293 (
            .O(N__45178),
            .I(N__45167));
    Span4Mux_v I__10292 (
            .O(N__45173),
            .I(N__45167));
    InMux I__10291 (
            .O(N__45172),
            .I(N__45164));
    Odrv4 I__10290 (
            .O(N__45167),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    LocalMux I__10289 (
            .O(N__45164),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    CascadeMux I__10288 (
            .O(N__45159),
            .I(N__45156));
    InMux I__10287 (
            .O(N__45156),
            .I(N__45153));
    LocalMux I__10286 (
            .O(N__45153),
            .I(N__45150));
    Odrv4 I__10285 (
            .O(N__45150),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    InMux I__10284 (
            .O(N__45147),
            .I(N__45143));
    InMux I__10283 (
            .O(N__45146),
            .I(N__45140));
    LocalMux I__10282 (
            .O(N__45143),
            .I(N__45136));
    LocalMux I__10281 (
            .O(N__45140),
            .I(N__45133));
    InMux I__10280 (
            .O(N__45139),
            .I(N__45130));
    Span4Mux_v I__10279 (
            .O(N__45136),
            .I(N__45127));
    Span4Mux_h I__10278 (
            .O(N__45133),
            .I(N__45124));
    LocalMux I__10277 (
            .O(N__45130),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__10276 (
            .O(N__45127),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__10275 (
            .O(N__45124),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__10274 (
            .O(N__45117),
            .I(N__45114));
    LocalMux I__10273 (
            .O(N__45114),
            .I(N__45111));
    Span4Mux_h I__10272 (
            .O(N__45111),
            .I(N__45108));
    Odrv4 I__10271 (
            .O(N__45108),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    InMux I__10270 (
            .O(N__45105),
            .I(N__45102));
    LocalMux I__10269 (
            .O(N__45102),
            .I(N__45099));
    Odrv4 I__10268 (
            .O(N__45099),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    InMux I__10267 (
            .O(N__45096),
            .I(N__45090));
    InMux I__10266 (
            .O(N__45095),
            .I(N__45090));
    LocalMux I__10265 (
            .O(N__45090),
            .I(N__45087));
    Odrv4 I__10264 (
            .O(N__45087),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__10263 (
            .O(N__45084),
            .I(N__45079));
    InMux I__10262 (
            .O(N__45083),
            .I(N__45076));
    InMux I__10261 (
            .O(N__45082),
            .I(N__45071));
    InMux I__10260 (
            .O(N__45079),
            .I(N__45071));
    LocalMux I__10259 (
            .O(N__45076),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__10258 (
            .O(N__45071),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__10257 (
            .O(N__45066),
            .I(N__45061));
    InMux I__10256 (
            .O(N__45065),
            .I(N__45056));
    InMux I__10255 (
            .O(N__45064),
            .I(N__45056));
    LocalMux I__10254 (
            .O(N__45061),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__10253 (
            .O(N__45056),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    CascadeMux I__10252 (
            .O(N__45051),
            .I(N__45048));
    InMux I__10251 (
            .O(N__45048),
            .I(N__45045));
    LocalMux I__10250 (
            .O(N__45045),
            .I(N__45042));
    Odrv12 I__10249 (
            .O(N__45042),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    InMux I__10248 (
            .O(N__45039),
            .I(N__45035));
    InMux I__10247 (
            .O(N__45038),
            .I(N__45031));
    LocalMux I__10246 (
            .O(N__45035),
            .I(N__45028));
    InMux I__10245 (
            .O(N__45034),
            .I(N__45025));
    LocalMux I__10244 (
            .O(N__45031),
            .I(N__45020));
    Span4Mux_v I__10243 (
            .O(N__45028),
            .I(N__45020));
    LocalMux I__10242 (
            .O(N__45025),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__10241 (
            .O(N__45020),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__10240 (
            .O(N__45015),
            .I(N__45010));
    InMux I__10239 (
            .O(N__45014),
            .I(N__45007));
    InMux I__10238 (
            .O(N__45013),
            .I(N__45004));
    LocalMux I__10237 (
            .O(N__45010),
            .I(N__45000));
    LocalMux I__10236 (
            .O(N__45007),
            .I(N__44997));
    LocalMux I__10235 (
            .O(N__45004),
            .I(N__44994));
    InMux I__10234 (
            .O(N__45003),
            .I(N__44991));
    Span4Mux_v I__10233 (
            .O(N__45000),
            .I(N__44988));
    Span12Mux_s11_v I__10232 (
            .O(N__44997),
            .I(N__44985));
    Span4Mux_v I__10231 (
            .O(N__44994),
            .I(N__44980));
    LocalMux I__10230 (
            .O(N__44991),
            .I(N__44980));
    Odrv4 I__10229 (
            .O(N__44988),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv12 I__10228 (
            .O(N__44985),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__10227 (
            .O(N__44980),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    CascadeMux I__10226 (
            .O(N__44973),
            .I(N__44969));
    InMux I__10225 (
            .O(N__44972),
            .I(N__44964));
    InMux I__10224 (
            .O(N__44969),
            .I(N__44964));
    LocalMux I__10223 (
            .O(N__44964),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    CascadeMux I__10222 (
            .O(N__44961),
            .I(N__44958));
    InMux I__10221 (
            .O(N__44958),
            .I(N__44955));
    LocalMux I__10220 (
            .O(N__44955),
            .I(N__44952));
    Odrv12 I__10219 (
            .O(N__44952),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    CascadeMux I__10218 (
            .O(N__44949),
            .I(N__44944));
    InMux I__10217 (
            .O(N__44948),
            .I(N__44941));
    InMux I__10216 (
            .O(N__44947),
            .I(N__44938));
    InMux I__10215 (
            .O(N__44944),
            .I(N__44935));
    LocalMux I__10214 (
            .O(N__44941),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__10213 (
            .O(N__44938),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__10212 (
            .O(N__44935),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__10211 (
            .O(N__44928),
            .I(N__44922));
    InMux I__10210 (
            .O(N__44927),
            .I(N__44922));
    LocalMux I__10209 (
            .O(N__44922),
            .I(N__44919));
    Odrv4 I__10208 (
            .O(N__44919),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    InMux I__10207 (
            .O(N__44916),
            .I(N__44911));
    InMux I__10206 (
            .O(N__44915),
            .I(N__44908));
    InMux I__10205 (
            .O(N__44914),
            .I(N__44905));
    LocalMux I__10204 (
            .O(N__44911),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__10203 (
            .O(N__44908),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__10202 (
            .O(N__44905),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__10201 (
            .O(N__44898),
            .I(N__44895));
    LocalMux I__10200 (
            .O(N__44895),
            .I(N__44892));
    Odrv4 I__10199 (
            .O(N__44892),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    InMux I__10198 (
            .O(N__44889),
            .I(N__44886));
    LocalMux I__10197 (
            .O(N__44886),
            .I(N__44883));
    Span4Mux_v I__10196 (
            .O(N__44883),
            .I(N__44880));
    Odrv4 I__10195 (
            .O(N__44880),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    InMux I__10194 (
            .O(N__44877),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__10193 (
            .O(N__44874),
            .I(N__44854));
    InMux I__10192 (
            .O(N__44873),
            .I(N__44854));
    InMux I__10191 (
            .O(N__44872),
            .I(N__44854));
    InMux I__10190 (
            .O(N__44871),
            .I(N__44854));
    InMux I__10189 (
            .O(N__44870),
            .I(N__44837));
    InMux I__10188 (
            .O(N__44869),
            .I(N__44837));
    InMux I__10187 (
            .O(N__44868),
            .I(N__44837));
    InMux I__10186 (
            .O(N__44867),
            .I(N__44837));
    InMux I__10185 (
            .O(N__44866),
            .I(N__44828));
    InMux I__10184 (
            .O(N__44865),
            .I(N__44828));
    InMux I__10183 (
            .O(N__44864),
            .I(N__44828));
    InMux I__10182 (
            .O(N__44863),
            .I(N__44828));
    LocalMux I__10181 (
            .O(N__44854),
            .I(N__44815));
    InMux I__10180 (
            .O(N__44853),
            .I(N__44806));
    InMux I__10179 (
            .O(N__44852),
            .I(N__44806));
    InMux I__10178 (
            .O(N__44851),
            .I(N__44806));
    InMux I__10177 (
            .O(N__44850),
            .I(N__44806));
    InMux I__10176 (
            .O(N__44849),
            .I(N__44797));
    InMux I__10175 (
            .O(N__44848),
            .I(N__44797));
    InMux I__10174 (
            .O(N__44847),
            .I(N__44797));
    InMux I__10173 (
            .O(N__44846),
            .I(N__44797));
    LocalMux I__10172 (
            .O(N__44837),
            .I(N__44792));
    LocalMux I__10171 (
            .O(N__44828),
            .I(N__44792));
    InMux I__10170 (
            .O(N__44827),
            .I(N__44787));
    InMux I__10169 (
            .O(N__44826),
            .I(N__44787));
    InMux I__10168 (
            .O(N__44825),
            .I(N__44778));
    InMux I__10167 (
            .O(N__44824),
            .I(N__44778));
    InMux I__10166 (
            .O(N__44823),
            .I(N__44778));
    InMux I__10165 (
            .O(N__44822),
            .I(N__44778));
    InMux I__10164 (
            .O(N__44821),
            .I(N__44769));
    InMux I__10163 (
            .O(N__44820),
            .I(N__44769));
    InMux I__10162 (
            .O(N__44819),
            .I(N__44769));
    InMux I__10161 (
            .O(N__44818),
            .I(N__44769));
    Span4Mux_v I__10160 (
            .O(N__44815),
            .I(N__44762));
    LocalMux I__10159 (
            .O(N__44806),
            .I(N__44762));
    LocalMux I__10158 (
            .O(N__44797),
            .I(N__44762));
    Span4Mux_v I__10157 (
            .O(N__44792),
            .I(N__44755));
    LocalMux I__10156 (
            .O(N__44787),
            .I(N__44755));
    LocalMux I__10155 (
            .O(N__44778),
            .I(N__44755));
    LocalMux I__10154 (
            .O(N__44769),
            .I(N__44752));
    Span4Mux_h I__10153 (
            .O(N__44762),
            .I(N__44749));
    Span4Mux_h I__10152 (
            .O(N__44755),
            .I(N__44746));
    Odrv12 I__10151 (
            .O(N__44752),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__10150 (
            .O(N__44749),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__10149 (
            .O(N__44746),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__10148 (
            .O(N__44739),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__10147 (
            .O(N__44736),
            .I(N__44733));
    InMux I__10146 (
            .O(N__44733),
            .I(N__44730));
    LocalMux I__10145 (
            .O(N__44730),
            .I(N__44726));
    InMux I__10144 (
            .O(N__44729),
            .I(N__44723));
    Span4Mux_h I__10143 (
            .O(N__44726),
            .I(N__44720));
    LocalMux I__10142 (
            .O(N__44723),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__10141 (
            .O(N__44720),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__10140 (
            .O(N__44715),
            .I(N__44710));
    CEMux I__10139 (
            .O(N__44714),
            .I(N__44707));
    CEMux I__10138 (
            .O(N__44713),
            .I(N__44703));
    LocalMux I__10137 (
            .O(N__44710),
            .I(N__44700));
    LocalMux I__10136 (
            .O(N__44707),
            .I(N__44697));
    CEMux I__10135 (
            .O(N__44706),
            .I(N__44694));
    LocalMux I__10134 (
            .O(N__44703),
            .I(N__44691));
    Span4Mux_v I__10133 (
            .O(N__44700),
            .I(N__44686));
    Span4Mux_h I__10132 (
            .O(N__44697),
            .I(N__44686));
    LocalMux I__10131 (
            .O(N__44694),
            .I(N__44683));
    Span4Mux_h I__10130 (
            .O(N__44691),
            .I(N__44680));
    Span4Mux_h I__10129 (
            .O(N__44686),
            .I(N__44677));
    Span4Mux_h I__10128 (
            .O(N__44683),
            .I(N__44674));
    Odrv4 I__10127 (
            .O(N__44680),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    Odrv4 I__10126 (
            .O(N__44677),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    Odrv4 I__10125 (
            .O(N__44674),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    InMux I__10124 (
            .O(N__44667),
            .I(N__44664));
    LocalMux I__10123 (
            .O(N__44664),
            .I(N__44658));
    InMux I__10122 (
            .O(N__44663),
            .I(N__44655));
    InMux I__10121 (
            .O(N__44662),
            .I(N__44650));
    InMux I__10120 (
            .O(N__44661),
            .I(N__44650));
    Span4Mux_v I__10119 (
            .O(N__44658),
            .I(N__44647));
    LocalMux I__10118 (
            .O(N__44655),
            .I(N__44644));
    LocalMux I__10117 (
            .O(N__44650),
            .I(N__44641));
    Span4Mux_v I__10116 (
            .O(N__44647),
            .I(N__44636));
    Span4Mux_v I__10115 (
            .O(N__44644),
            .I(N__44636));
    Odrv4 I__10114 (
            .O(N__44641),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__10113 (
            .O(N__44636),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__10112 (
            .O(N__44631),
            .I(N__44628));
    LocalMux I__10111 (
            .O(N__44628),
            .I(N__44625));
    Span4Mux_h I__10110 (
            .O(N__44625),
            .I(N__44621));
    InMux I__10109 (
            .O(N__44624),
            .I(N__44618));
    Odrv4 I__10108 (
            .O(N__44621),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__10107 (
            .O(N__44618),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    InMux I__10106 (
            .O(N__44613),
            .I(N__44608));
    InMux I__10105 (
            .O(N__44612),
            .I(N__44605));
    InMux I__10104 (
            .O(N__44611),
            .I(N__44602));
    LocalMux I__10103 (
            .O(N__44608),
            .I(N__44599));
    LocalMux I__10102 (
            .O(N__44605),
            .I(N__44596));
    LocalMux I__10101 (
            .O(N__44602),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    Odrv4 I__10100 (
            .O(N__44599),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    Odrv4 I__10099 (
            .O(N__44596),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    InMux I__10098 (
            .O(N__44589),
            .I(N__44585));
    InMux I__10097 (
            .O(N__44588),
            .I(N__44581));
    LocalMux I__10096 (
            .O(N__44585),
            .I(N__44578));
    InMux I__10095 (
            .O(N__44584),
            .I(N__44575));
    LocalMux I__10094 (
            .O(N__44581),
            .I(N__44571));
    Span4Mux_v I__10093 (
            .O(N__44578),
            .I(N__44566));
    LocalMux I__10092 (
            .O(N__44575),
            .I(N__44566));
    InMux I__10091 (
            .O(N__44574),
            .I(N__44563));
    Span12Mux_s10_v I__10090 (
            .O(N__44571),
            .I(N__44560));
    Span4Mux_v I__10089 (
            .O(N__44566),
            .I(N__44557));
    LocalMux I__10088 (
            .O(N__44563),
            .I(N__44554));
    Odrv12 I__10087 (
            .O(N__44560),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__10086 (
            .O(N__44557),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__10085 (
            .O(N__44554),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__10084 (
            .O(N__44547),
            .I(N__44542));
    InMux I__10083 (
            .O(N__44546),
            .I(N__44537));
    InMux I__10082 (
            .O(N__44545),
            .I(N__44537));
    LocalMux I__10081 (
            .O(N__44542),
            .I(N__44534));
    LocalMux I__10080 (
            .O(N__44537),
            .I(N__44531));
    Span4Mux_h I__10079 (
            .O(N__44534),
            .I(N__44525));
    Span4Mux_h I__10078 (
            .O(N__44531),
            .I(N__44525));
    InMux I__10077 (
            .O(N__44530),
            .I(N__44522));
    Odrv4 I__10076 (
            .O(N__44525),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    LocalMux I__10075 (
            .O(N__44522),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__10074 (
            .O(N__44517),
            .I(N__44514));
    LocalMux I__10073 (
            .O(N__44514),
            .I(N__44510));
    InMux I__10072 (
            .O(N__44513),
            .I(N__44507));
    Odrv4 I__10071 (
            .O(N__44510),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    LocalMux I__10070 (
            .O(N__44507),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    InMux I__10069 (
            .O(N__44502),
            .I(N__44499));
    LocalMux I__10068 (
            .O(N__44499),
            .I(N__44496));
    Span4Mux_h I__10067 (
            .O(N__44496),
            .I(N__44493));
    Odrv4 I__10066 (
            .O(N__44493),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    InMux I__10065 (
            .O(N__44490),
            .I(N__44487));
    LocalMux I__10064 (
            .O(N__44487),
            .I(N__44484));
    Span4Mux_v I__10063 (
            .O(N__44484),
            .I(N__44481));
    Odrv4 I__10062 (
            .O(N__44481),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    CascadeMux I__10061 (
            .O(N__44478),
            .I(N__44473));
    InMux I__10060 (
            .O(N__44477),
            .I(N__44470));
    InMux I__10059 (
            .O(N__44476),
            .I(N__44465));
    InMux I__10058 (
            .O(N__44473),
            .I(N__44465));
    LocalMux I__10057 (
            .O(N__44470),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__10056 (
            .O(N__44465),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__10055 (
            .O(N__44460),
            .I(N__44455));
    InMux I__10054 (
            .O(N__44459),
            .I(N__44452));
    InMux I__10053 (
            .O(N__44458),
            .I(N__44447));
    InMux I__10052 (
            .O(N__44455),
            .I(N__44447));
    LocalMux I__10051 (
            .O(N__44452),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__10050 (
            .O(N__44447),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__10049 (
            .O(N__44442),
            .I(N__44436));
    InMux I__10048 (
            .O(N__44441),
            .I(N__44436));
    LocalMux I__10047 (
            .O(N__44436),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__10046 (
            .O(N__44433),
            .I(N__44430));
    InMux I__10045 (
            .O(N__44430),
            .I(N__44427));
    LocalMux I__10044 (
            .O(N__44427),
            .I(N__44424));
    Span4Mux_h I__10043 (
            .O(N__44424),
            .I(N__44421));
    Odrv4 I__10042 (
            .O(N__44421),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    InMux I__10041 (
            .O(N__44418),
            .I(N__44413));
    InMux I__10040 (
            .O(N__44417),
            .I(N__44408));
    InMux I__10039 (
            .O(N__44416),
            .I(N__44408));
    LocalMux I__10038 (
            .O(N__44413),
            .I(N__44404));
    LocalMux I__10037 (
            .O(N__44408),
            .I(N__44401));
    CascadeMux I__10036 (
            .O(N__44407),
            .I(N__44398));
    Span4Mux_v I__10035 (
            .O(N__44404),
            .I(N__44395));
    Span4Mux_h I__10034 (
            .O(N__44401),
            .I(N__44392));
    InMux I__10033 (
            .O(N__44398),
            .I(N__44389));
    Odrv4 I__10032 (
            .O(N__44395),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__10031 (
            .O(N__44392),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__10030 (
            .O(N__44389),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__10029 (
            .O(N__44382),
            .I(N__44379));
    LocalMux I__10028 (
            .O(N__44379),
            .I(N__44376));
    Span4Mux_h I__10027 (
            .O(N__44376),
            .I(N__44372));
    InMux I__10026 (
            .O(N__44375),
            .I(N__44369));
    Odrv4 I__10025 (
            .O(N__44372),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    LocalMux I__10024 (
            .O(N__44369),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__10023 (
            .O(N__44364),
            .I(N__44358));
    InMux I__10022 (
            .O(N__44363),
            .I(N__44358));
    LocalMux I__10021 (
            .O(N__44358),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__10020 (
            .O(N__44355),
            .I(N__44351));
    InMux I__10019 (
            .O(N__44354),
            .I(N__44348));
    LocalMux I__10018 (
            .O(N__44351),
            .I(N__44344));
    LocalMux I__10017 (
            .O(N__44348),
            .I(N__44341));
    InMux I__10016 (
            .O(N__44347),
            .I(N__44338));
    Span4Mux_v I__10015 (
            .O(N__44344),
            .I(N__44335));
    Span4Mux_v I__10014 (
            .O(N__44341),
            .I(N__44332));
    LocalMux I__10013 (
            .O(N__44338),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    Odrv4 I__10012 (
            .O(N__44335),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    Odrv4 I__10011 (
            .O(N__44332),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    InMux I__10010 (
            .O(N__44325),
            .I(N__44322));
    LocalMux I__10009 (
            .O(N__44322),
            .I(N__44317));
    InMux I__10008 (
            .O(N__44321),
            .I(N__44314));
    InMux I__10007 (
            .O(N__44320),
            .I(N__44311));
    Span4Mux_h I__10006 (
            .O(N__44317),
            .I(N__44307));
    LocalMux I__10005 (
            .O(N__44314),
            .I(N__44304));
    LocalMux I__10004 (
            .O(N__44311),
            .I(N__44301));
    InMux I__10003 (
            .O(N__44310),
            .I(N__44298));
    Odrv4 I__10002 (
            .O(N__44307),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv12 I__10001 (
            .O(N__44304),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__10000 (
            .O(N__44301),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__9999 (
            .O(N__44298),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    CascadeMux I__9998 (
            .O(N__44289),
            .I(N__44285));
    CascadeMux I__9997 (
            .O(N__44288),
            .I(N__44282));
    InMux I__9996 (
            .O(N__44285),
            .I(N__44277));
    InMux I__9995 (
            .O(N__44282),
            .I(N__44277));
    LocalMux I__9994 (
            .O(N__44277),
            .I(N__44273));
    InMux I__9993 (
            .O(N__44276),
            .I(N__44270));
    Span4Mux_h I__9992 (
            .O(N__44273),
            .I(N__44267));
    LocalMux I__9991 (
            .O(N__44270),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__9990 (
            .O(N__44267),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__9989 (
            .O(N__44262),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__9988 (
            .O(N__44259),
            .I(N__44255));
    CascadeMux I__9987 (
            .O(N__44258),
            .I(N__44252));
    InMux I__9986 (
            .O(N__44255),
            .I(N__44247));
    InMux I__9985 (
            .O(N__44252),
            .I(N__44247));
    LocalMux I__9984 (
            .O(N__44247),
            .I(N__44243));
    InMux I__9983 (
            .O(N__44246),
            .I(N__44240));
    Span4Mux_v I__9982 (
            .O(N__44243),
            .I(N__44237));
    LocalMux I__9981 (
            .O(N__44240),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__9980 (
            .O(N__44237),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__9979 (
            .O(N__44232),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__9978 (
            .O(N__44229),
            .I(N__44223));
    InMux I__9977 (
            .O(N__44228),
            .I(N__44223));
    LocalMux I__9976 (
            .O(N__44223),
            .I(N__44219));
    InMux I__9975 (
            .O(N__44222),
            .I(N__44216));
    Span4Mux_v I__9974 (
            .O(N__44219),
            .I(N__44213));
    LocalMux I__9973 (
            .O(N__44216),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__9972 (
            .O(N__44213),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__9971 (
            .O(N__44208),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__9970 (
            .O(N__44205),
            .I(N__44202));
    InMux I__9969 (
            .O(N__44202),
            .I(N__44198));
    InMux I__9968 (
            .O(N__44201),
            .I(N__44195));
    LocalMux I__9967 (
            .O(N__44198),
            .I(N__44189));
    LocalMux I__9966 (
            .O(N__44195),
            .I(N__44189));
    InMux I__9965 (
            .O(N__44194),
            .I(N__44186));
    Span4Mux_v I__9964 (
            .O(N__44189),
            .I(N__44183));
    LocalMux I__9963 (
            .O(N__44186),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__9962 (
            .O(N__44183),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__9961 (
            .O(N__44178),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__9960 (
            .O(N__44175),
            .I(N__44171));
    CascadeMux I__9959 (
            .O(N__44174),
            .I(N__44168));
    InMux I__9958 (
            .O(N__44171),
            .I(N__44165));
    InMux I__9957 (
            .O(N__44168),
            .I(N__44162));
    LocalMux I__9956 (
            .O(N__44165),
            .I(N__44156));
    LocalMux I__9955 (
            .O(N__44162),
            .I(N__44156));
    InMux I__9954 (
            .O(N__44161),
            .I(N__44153));
    Sp12to4 I__9953 (
            .O(N__44156),
            .I(N__44150));
    LocalMux I__9952 (
            .O(N__44153),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv12 I__9951 (
            .O(N__44150),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__9950 (
            .O(N__44145),
            .I(bfn_17_26_0_));
    CascadeMux I__9949 (
            .O(N__44142),
            .I(N__44139));
    InMux I__9948 (
            .O(N__44139),
            .I(N__44135));
    InMux I__9947 (
            .O(N__44138),
            .I(N__44132));
    LocalMux I__9946 (
            .O(N__44135),
            .I(N__44128));
    LocalMux I__9945 (
            .O(N__44132),
            .I(N__44125));
    InMux I__9944 (
            .O(N__44131),
            .I(N__44122));
    Span4Mux_h I__9943 (
            .O(N__44128),
            .I(N__44119));
    Span4Mux_v I__9942 (
            .O(N__44125),
            .I(N__44116));
    LocalMux I__9941 (
            .O(N__44122),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__9940 (
            .O(N__44119),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__9939 (
            .O(N__44116),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__9938 (
            .O(N__44109),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__9937 (
            .O(N__44106),
            .I(N__44103));
    InMux I__9936 (
            .O(N__44103),
            .I(N__44099));
    InMux I__9935 (
            .O(N__44102),
            .I(N__44096));
    LocalMux I__9934 (
            .O(N__44099),
            .I(N__44090));
    LocalMux I__9933 (
            .O(N__44096),
            .I(N__44090));
    InMux I__9932 (
            .O(N__44095),
            .I(N__44087));
    Span4Mux_h I__9931 (
            .O(N__44090),
            .I(N__44084));
    LocalMux I__9930 (
            .O(N__44087),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__9929 (
            .O(N__44084),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__9928 (
            .O(N__44079),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__9927 (
            .O(N__44076),
            .I(N__44070));
    InMux I__9926 (
            .O(N__44075),
            .I(N__44070));
    LocalMux I__9925 (
            .O(N__44070),
            .I(N__44066));
    InMux I__9924 (
            .O(N__44069),
            .I(N__44063));
    Span4Mux_h I__9923 (
            .O(N__44066),
            .I(N__44060));
    LocalMux I__9922 (
            .O(N__44063),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__9921 (
            .O(N__44060),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__9920 (
            .O(N__44055),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__9919 (
            .O(N__44052),
            .I(N__44049));
    LocalMux I__9918 (
            .O(N__44049),
            .I(N__44045));
    InMux I__9917 (
            .O(N__44048),
            .I(N__44042));
    Span4Mux_h I__9916 (
            .O(N__44045),
            .I(N__44039));
    LocalMux I__9915 (
            .O(N__44042),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__9914 (
            .O(N__44039),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__9913 (
            .O(N__44034),
            .I(N__44028));
    InMux I__9912 (
            .O(N__44033),
            .I(N__44028));
    LocalMux I__9911 (
            .O(N__44028),
            .I(N__44024));
    InMux I__9910 (
            .O(N__44027),
            .I(N__44021));
    Span4Mux_h I__9909 (
            .O(N__44024),
            .I(N__44018));
    LocalMux I__9908 (
            .O(N__44021),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__9907 (
            .O(N__44018),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__9906 (
            .O(N__44013),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__9905 (
            .O(N__44010),
            .I(N__44006));
    CascadeMux I__9904 (
            .O(N__44009),
            .I(N__44003));
    InMux I__9903 (
            .O(N__44006),
            .I(N__43998));
    InMux I__9902 (
            .O(N__44003),
            .I(N__43998));
    LocalMux I__9901 (
            .O(N__43998),
            .I(N__43994));
    InMux I__9900 (
            .O(N__43997),
            .I(N__43991));
    Span4Mux_h I__9899 (
            .O(N__43994),
            .I(N__43988));
    LocalMux I__9898 (
            .O(N__43991),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__9897 (
            .O(N__43988),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__9896 (
            .O(N__43983),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__9895 (
            .O(N__43980),
            .I(N__43976));
    CascadeMux I__9894 (
            .O(N__43979),
            .I(N__43973));
    InMux I__9893 (
            .O(N__43976),
            .I(N__43968));
    InMux I__9892 (
            .O(N__43973),
            .I(N__43968));
    LocalMux I__9891 (
            .O(N__43968),
            .I(N__43964));
    InMux I__9890 (
            .O(N__43967),
            .I(N__43961));
    Span4Mux_v I__9889 (
            .O(N__43964),
            .I(N__43958));
    LocalMux I__9888 (
            .O(N__43961),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__9887 (
            .O(N__43958),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__9886 (
            .O(N__43953),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    CascadeMux I__9885 (
            .O(N__43950),
            .I(N__43947));
    InMux I__9884 (
            .O(N__43947),
            .I(N__43943));
    InMux I__9883 (
            .O(N__43946),
            .I(N__43940));
    LocalMux I__9882 (
            .O(N__43943),
            .I(N__43934));
    LocalMux I__9881 (
            .O(N__43940),
            .I(N__43934));
    InMux I__9880 (
            .O(N__43939),
            .I(N__43931));
    Span4Mux_v I__9879 (
            .O(N__43934),
            .I(N__43928));
    LocalMux I__9878 (
            .O(N__43931),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__9877 (
            .O(N__43928),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__9876 (
            .O(N__43923),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__9875 (
            .O(N__43920),
            .I(N__43917));
    InMux I__9874 (
            .O(N__43917),
            .I(N__43913));
    InMux I__9873 (
            .O(N__43916),
            .I(N__43910));
    LocalMux I__9872 (
            .O(N__43913),
            .I(N__43904));
    LocalMux I__9871 (
            .O(N__43910),
            .I(N__43904));
    InMux I__9870 (
            .O(N__43909),
            .I(N__43901));
    Span4Mux_v I__9869 (
            .O(N__43904),
            .I(N__43898));
    LocalMux I__9868 (
            .O(N__43901),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__9867 (
            .O(N__43898),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__9866 (
            .O(N__43893),
            .I(bfn_17_25_0_));
    CascadeMux I__9865 (
            .O(N__43890),
            .I(N__43887));
    InMux I__9864 (
            .O(N__43887),
            .I(N__43883));
    InMux I__9863 (
            .O(N__43886),
            .I(N__43880));
    LocalMux I__9862 (
            .O(N__43883),
            .I(N__43876));
    LocalMux I__9861 (
            .O(N__43880),
            .I(N__43873));
    InMux I__9860 (
            .O(N__43879),
            .I(N__43870));
    Span4Mux_h I__9859 (
            .O(N__43876),
            .I(N__43867));
    Span4Mux_v I__9858 (
            .O(N__43873),
            .I(N__43864));
    LocalMux I__9857 (
            .O(N__43870),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__9856 (
            .O(N__43867),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__9855 (
            .O(N__43864),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__9854 (
            .O(N__43857),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__9853 (
            .O(N__43854),
            .I(N__43848));
    InMux I__9852 (
            .O(N__43853),
            .I(N__43848));
    LocalMux I__9851 (
            .O(N__43848),
            .I(N__43844));
    InMux I__9850 (
            .O(N__43847),
            .I(N__43841));
    Span4Mux_h I__9849 (
            .O(N__43844),
            .I(N__43838));
    LocalMux I__9848 (
            .O(N__43841),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__9847 (
            .O(N__43838),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__9846 (
            .O(N__43833),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__9845 (
            .O(N__43830),
            .I(N__43824));
    InMux I__9844 (
            .O(N__43829),
            .I(N__43824));
    LocalMux I__9843 (
            .O(N__43824),
            .I(N__43820));
    InMux I__9842 (
            .O(N__43823),
            .I(N__43817));
    Span4Mux_h I__9841 (
            .O(N__43820),
            .I(N__43814));
    LocalMux I__9840 (
            .O(N__43817),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__9839 (
            .O(N__43814),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__9838 (
            .O(N__43809),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__9837 (
            .O(N__43806),
            .I(N__43802));
    CascadeMux I__9836 (
            .O(N__43805),
            .I(N__43799));
    InMux I__9835 (
            .O(N__43802),
            .I(N__43794));
    InMux I__9834 (
            .O(N__43799),
            .I(N__43794));
    LocalMux I__9833 (
            .O(N__43794),
            .I(N__43790));
    InMux I__9832 (
            .O(N__43793),
            .I(N__43787));
    Span4Mux_h I__9831 (
            .O(N__43790),
            .I(N__43784));
    LocalMux I__9830 (
            .O(N__43787),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__9829 (
            .O(N__43784),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__9828 (
            .O(N__43779),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__9827 (
            .O(N__43776),
            .I(N__43772));
    CascadeMux I__9826 (
            .O(N__43775),
            .I(N__43769));
    InMux I__9825 (
            .O(N__43772),
            .I(N__43764));
    InMux I__9824 (
            .O(N__43769),
            .I(N__43764));
    LocalMux I__9823 (
            .O(N__43764),
            .I(N__43760));
    InMux I__9822 (
            .O(N__43763),
            .I(N__43757));
    Span4Mux_v I__9821 (
            .O(N__43760),
            .I(N__43754));
    LocalMux I__9820 (
            .O(N__43757),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__9819 (
            .O(N__43754),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__9818 (
            .O(N__43749),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__9817 (
            .O(N__43746),
            .I(N__43743));
    InMux I__9816 (
            .O(N__43743),
            .I(N__43739));
    InMux I__9815 (
            .O(N__43742),
            .I(N__43736));
    LocalMux I__9814 (
            .O(N__43739),
            .I(N__43730));
    LocalMux I__9813 (
            .O(N__43736),
            .I(N__43730));
    InMux I__9812 (
            .O(N__43735),
            .I(N__43727));
    Span4Mux_h I__9811 (
            .O(N__43730),
            .I(N__43724));
    LocalMux I__9810 (
            .O(N__43727),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__9809 (
            .O(N__43724),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__9808 (
            .O(N__43719),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__9807 (
            .O(N__43716),
            .I(N__43710));
    InMux I__9806 (
            .O(N__43715),
            .I(N__43710));
    LocalMux I__9805 (
            .O(N__43710),
            .I(N__43706));
    InMux I__9804 (
            .O(N__43709),
            .I(N__43703));
    Span4Mux_v I__9803 (
            .O(N__43706),
            .I(N__43700));
    LocalMux I__9802 (
            .O(N__43703),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__9801 (
            .O(N__43700),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__9800 (
            .O(N__43695),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__9799 (
            .O(N__43692),
            .I(N__43686));
    InMux I__9798 (
            .O(N__43691),
            .I(N__43686));
    LocalMux I__9797 (
            .O(N__43686),
            .I(N__43682));
    InMux I__9796 (
            .O(N__43685),
            .I(N__43679));
    Span4Mux_v I__9795 (
            .O(N__43682),
            .I(N__43676));
    LocalMux I__9794 (
            .O(N__43679),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__9793 (
            .O(N__43676),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__9792 (
            .O(N__43671),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__9791 (
            .O(N__43668),
            .I(N__43664));
    CascadeMux I__9790 (
            .O(N__43667),
            .I(N__43661));
    InMux I__9789 (
            .O(N__43664),
            .I(N__43658));
    InMux I__9788 (
            .O(N__43661),
            .I(N__43655));
    LocalMux I__9787 (
            .O(N__43658),
            .I(N__43649));
    LocalMux I__9786 (
            .O(N__43655),
            .I(N__43649));
    InMux I__9785 (
            .O(N__43654),
            .I(N__43646));
    Span4Mux_v I__9784 (
            .O(N__43649),
            .I(N__43643));
    LocalMux I__9783 (
            .O(N__43646),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__9782 (
            .O(N__43643),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__9781 (
            .O(N__43638),
            .I(bfn_17_24_0_));
    CascadeMux I__9780 (
            .O(N__43635),
            .I(N__43631));
    CascadeMux I__9779 (
            .O(N__43634),
            .I(N__43628));
    InMux I__9778 (
            .O(N__43631),
            .I(N__43625));
    InMux I__9777 (
            .O(N__43628),
            .I(N__43622));
    LocalMux I__9776 (
            .O(N__43625),
            .I(N__43619));
    LocalMux I__9775 (
            .O(N__43622),
            .I(N__43615));
    Span4Mux_v I__9774 (
            .O(N__43619),
            .I(N__43612));
    InMux I__9773 (
            .O(N__43618),
            .I(N__43609));
    Span4Mux_h I__9772 (
            .O(N__43615),
            .I(N__43604));
    Span4Mux_h I__9771 (
            .O(N__43612),
            .I(N__43604));
    LocalMux I__9770 (
            .O(N__43609),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__9769 (
            .O(N__43604),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__9768 (
            .O(N__43599),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__9767 (
            .O(N__43596),
            .I(N__43593));
    InMux I__9766 (
            .O(N__43593),
            .I(N__43589));
    InMux I__9765 (
            .O(N__43592),
            .I(N__43586));
    LocalMux I__9764 (
            .O(N__43589),
            .I(N__43580));
    LocalMux I__9763 (
            .O(N__43586),
            .I(N__43580));
    InMux I__9762 (
            .O(N__43585),
            .I(N__43577));
    Span4Mux_h I__9761 (
            .O(N__43580),
            .I(N__43574));
    LocalMux I__9760 (
            .O(N__43577),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__9759 (
            .O(N__43574),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__9758 (
            .O(N__43569),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__9757 (
            .O(N__43566),
            .I(N__43560));
    InMux I__9756 (
            .O(N__43565),
            .I(N__43560));
    LocalMux I__9755 (
            .O(N__43560),
            .I(N__43556));
    InMux I__9754 (
            .O(N__43559),
            .I(N__43553));
    Span4Mux_h I__9753 (
            .O(N__43556),
            .I(N__43550));
    LocalMux I__9752 (
            .O(N__43553),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__9751 (
            .O(N__43550),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__9750 (
            .O(N__43545),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__9749 (
            .O(N__43542),
            .I(N__43539));
    LocalMux I__9748 (
            .O(N__43539),
            .I(N__43536));
    Odrv12 I__9747 (
            .O(N__43536),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    CascadeMux I__9746 (
            .O(N__43533),
            .I(N__43529));
    CascadeMux I__9745 (
            .O(N__43532),
            .I(N__43526));
    InMux I__9744 (
            .O(N__43529),
            .I(N__43523));
    InMux I__9743 (
            .O(N__43526),
            .I(N__43520));
    LocalMux I__9742 (
            .O(N__43523),
            .I(N__43514));
    LocalMux I__9741 (
            .O(N__43520),
            .I(N__43514));
    InMux I__9740 (
            .O(N__43519),
            .I(N__43511));
    Span4Mux_h I__9739 (
            .O(N__43514),
            .I(N__43507));
    LocalMux I__9738 (
            .O(N__43511),
            .I(N__43504));
    InMux I__9737 (
            .O(N__43510),
            .I(N__43501));
    Odrv4 I__9736 (
            .O(N__43507),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__9735 (
            .O(N__43504),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__9734 (
            .O(N__43501),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__9733 (
            .O(N__43494),
            .I(N__43491));
    LocalMux I__9732 (
            .O(N__43491),
            .I(N__43488));
    Odrv12 I__9731 (
            .O(N__43488),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__9730 (
            .O(N__43485),
            .I(N__43481));
    InMux I__9729 (
            .O(N__43484),
            .I(N__43477));
    LocalMux I__9728 (
            .O(N__43481),
            .I(N__43474));
    InMux I__9727 (
            .O(N__43480),
            .I(N__43471));
    LocalMux I__9726 (
            .O(N__43477),
            .I(N__43465));
    Span4Mux_v I__9725 (
            .O(N__43474),
            .I(N__43465));
    LocalMux I__9724 (
            .O(N__43471),
            .I(N__43462));
    InMux I__9723 (
            .O(N__43470),
            .I(N__43459));
    Odrv4 I__9722 (
            .O(N__43465),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__9721 (
            .O(N__43462),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__9720 (
            .O(N__43459),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    CascadeMux I__9719 (
            .O(N__43452),
            .I(N__43449));
    InMux I__9718 (
            .O(N__43449),
            .I(N__43445));
    CascadeMux I__9717 (
            .O(N__43448),
            .I(N__43442));
    LocalMux I__9716 (
            .O(N__43445),
            .I(N__43438));
    InMux I__9715 (
            .O(N__43442),
            .I(N__43435));
    InMux I__9714 (
            .O(N__43441),
            .I(N__43432));
    Span4Mux_v I__9713 (
            .O(N__43438),
            .I(N__43429));
    LocalMux I__9712 (
            .O(N__43435),
            .I(N__43426));
    LocalMux I__9711 (
            .O(N__43432),
            .I(N__43423));
    Span4Mux_h I__9710 (
            .O(N__43429),
            .I(N__43420));
    Span4Mux_h I__9709 (
            .O(N__43426),
            .I(N__43417));
    Span4Mux_v I__9708 (
            .O(N__43423),
            .I(N__43414));
    Odrv4 I__9707 (
            .O(N__43420),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__9706 (
            .O(N__43417),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__9705 (
            .O(N__43414),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__9704 (
            .O(N__43407),
            .I(N__43404));
    InMux I__9703 (
            .O(N__43404),
            .I(N__43401));
    LocalMux I__9702 (
            .O(N__43401),
            .I(N__43398));
    Span4Mux_h I__9701 (
            .O(N__43398),
            .I(N__43395));
    Odrv4 I__9700 (
            .O(N__43395),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__9699 (
            .O(N__43392),
            .I(N__43389));
    LocalMux I__9698 (
            .O(N__43389),
            .I(N__43386));
    Odrv4 I__9697 (
            .O(N__43386),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__9696 (
            .O(N__43383),
            .I(N__43379));
    InMux I__9695 (
            .O(N__43382),
            .I(N__43376));
    InMux I__9694 (
            .O(N__43379),
            .I(N__43372));
    LocalMux I__9693 (
            .O(N__43376),
            .I(N__43368));
    InMux I__9692 (
            .O(N__43375),
            .I(N__43365));
    LocalMux I__9691 (
            .O(N__43372),
            .I(N__43362));
    InMux I__9690 (
            .O(N__43371),
            .I(N__43359));
    Span4Mux_h I__9689 (
            .O(N__43368),
            .I(N__43354));
    LocalMux I__9688 (
            .O(N__43365),
            .I(N__43354));
    Span4Mux_v I__9687 (
            .O(N__43362),
            .I(N__43349));
    LocalMux I__9686 (
            .O(N__43359),
            .I(N__43349));
    Odrv4 I__9685 (
            .O(N__43354),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__9684 (
            .O(N__43349),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__9683 (
            .O(N__43344),
            .I(N__43340));
    InMux I__9682 (
            .O(N__43343),
            .I(N__43337));
    LocalMux I__9681 (
            .O(N__43340),
            .I(N__43333));
    LocalMux I__9680 (
            .O(N__43337),
            .I(N__43330));
    InMux I__9679 (
            .O(N__43336),
            .I(N__43327));
    Span12Mux_h I__9678 (
            .O(N__43333),
            .I(N__43324));
    Span12Mux_h I__9677 (
            .O(N__43330),
            .I(N__43319));
    LocalMux I__9676 (
            .O(N__43327),
            .I(N__43319));
    Odrv12 I__9675 (
            .O(N__43324),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv12 I__9674 (
            .O(N__43319),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__9673 (
            .O(N__43314),
            .I(N__43311));
    LocalMux I__9672 (
            .O(N__43311),
            .I(N__43308));
    Odrv12 I__9671 (
            .O(N__43308),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__9670 (
            .O(N__43305),
            .I(bfn_17_23_0_));
    InMux I__9669 (
            .O(N__43302),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__9668 (
            .O(N__43299),
            .I(N__43295));
    InMux I__9667 (
            .O(N__43298),
            .I(N__43292));
    InMux I__9666 (
            .O(N__43295),
            .I(N__43289));
    LocalMux I__9665 (
            .O(N__43292),
            .I(N__43283));
    LocalMux I__9664 (
            .O(N__43289),
            .I(N__43283));
    InMux I__9663 (
            .O(N__43288),
            .I(N__43280));
    Sp12to4 I__9662 (
            .O(N__43283),
            .I(N__43277));
    LocalMux I__9661 (
            .O(N__43280),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__9660 (
            .O(N__43277),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__9659 (
            .O(N__43272),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__9658 (
            .O(N__43269),
            .I(N__43266));
    LocalMux I__9657 (
            .O(N__43266),
            .I(N__43263));
    Odrv12 I__9656 (
            .O(N__43263),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    CascadeMux I__9655 (
            .O(N__43260),
            .I(N__43257));
    InMux I__9654 (
            .O(N__43257),
            .I(N__43253));
    InMux I__9653 (
            .O(N__43256),
            .I(N__43250));
    LocalMux I__9652 (
            .O(N__43253),
            .I(N__43246));
    LocalMux I__9651 (
            .O(N__43250),
            .I(N__43243));
    InMux I__9650 (
            .O(N__43249),
            .I(N__43240));
    Span4Mux_h I__9649 (
            .O(N__43246),
            .I(N__43236));
    Span4Mux_v I__9648 (
            .O(N__43243),
            .I(N__43233));
    LocalMux I__9647 (
            .O(N__43240),
            .I(N__43230));
    InMux I__9646 (
            .O(N__43239),
            .I(N__43227));
    Odrv4 I__9645 (
            .O(N__43236),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__9644 (
            .O(N__43233),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv12 I__9643 (
            .O(N__43230),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__9642 (
            .O(N__43227),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__9641 (
            .O(N__43218),
            .I(N__43215));
    LocalMux I__9640 (
            .O(N__43215),
            .I(N__43212));
    Odrv12 I__9639 (
            .O(N__43212),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    CascadeMux I__9638 (
            .O(N__43209),
            .I(N__43206));
    InMux I__9637 (
            .O(N__43206),
            .I(N__43202));
    InMux I__9636 (
            .O(N__43205),
            .I(N__43198));
    LocalMux I__9635 (
            .O(N__43202),
            .I(N__43195));
    InMux I__9634 (
            .O(N__43201),
            .I(N__43192));
    LocalMux I__9633 (
            .O(N__43198),
            .I(N__43188));
    Span4Mux_v I__9632 (
            .O(N__43195),
            .I(N__43183));
    LocalMux I__9631 (
            .O(N__43192),
            .I(N__43183));
    InMux I__9630 (
            .O(N__43191),
            .I(N__43180));
    Odrv4 I__9629 (
            .O(N__43188),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__9628 (
            .O(N__43183),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__9627 (
            .O(N__43180),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__9626 (
            .O(N__43173),
            .I(N__43170));
    LocalMux I__9625 (
            .O(N__43170),
            .I(N__43167));
    Odrv4 I__9624 (
            .O(N__43167),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__9623 (
            .O(N__43164),
            .I(N__43160));
    CascadeMux I__9622 (
            .O(N__43163),
            .I(N__43157));
    LocalMux I__9621 (
            .O(N__43160),
            .I(N__43154));
    InMux I__9620 (
            .O(N__43157),
            .I(N__43151));
    Span4Mux_h I__9619 (
            .O(N__43154),
            .I(N__43147));
    LocalMux I__9618 (
            .O(N__43151),
            .I(N__43144));
    InMux I__9617 (
            .O(N__43150),
            .I(N__43141));
    Span4Mux_h I__9616 (
            .O(N__43147),
            .I(N__43135));
    Span4Mux_v I__9615 (
            .O(N__43144),
            .I(N__43135));
    LocalMux I__9614 (
            .O(N__43141),
            .I(N__43132));
    InMux I__9613 (
            .O(N__43140),
            .I(N__43129));
    Odrv4 I__9612 (
            .O(N__43135),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__9611 (
            .O(N__43132),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__9610 (
            .O(N__43129),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    CascadeMux I__9609 (
            .O(N__43122),
            .I(N__43119));
    InMux I__9608 (
            .O(N__43119),
            .I(N__43116));
    LocalMux I__9607 (
            .O(N__43116),
            .I(N__43113));
    Odrv4 I__9606 (
            .O(N__43113),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    CascadeMux I__9605 (
            .O(N__43110),
            .I(N__43107));
    InMux I__9604 (
            .O(N__43107),
            .I(N__43104));
    LocalMux I__9603 (
            .O(N__43104),
            .I(N__43099));
    InMux I__9602 (
            .O(N__43103),
            .I(N__43096));
    InMux I__9601 (
            .O(N__43102),
            .I(N__43093));
    Span12Mux_v I__9600 (
            .O(N__43099),
            .I(N__43089));
    LocalMux I__9599 (
            .O(N__43096),
            .I(N__43084));
    LocalMux I__9598 (
            .O(N__43093),
            .I(N__43084));
    InMux I__9597 (
            .O(N__43092),
            .I(N__43081));
    Odrv12 I__9596 (
            .O(N__43089),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv12 I__9595 (
            .O(N__43084),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__9594 (
            .O(N__43081),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__9593 (
            .O(N__43074),
            .I(N__43071));
    LocalMux I__9592 (
            .O(N__43071),
            .I(N__43068));
    Span4Mux_v I__9591 (
            .O(N__43068),
            .I(N__43065));
    Odrv4 I__9590 (
            .O(N__43065),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    CascadeMux I__9589 (
            .O(N__43062),
            .I(N__43058));
    CascadeMux I__9588 (
            .O(N__43061),
            .I(N__43055));
    InMux I__9587 (
            .O(N__43058),
            .I(N__43052));
    InMux I__9586 (
            .O(N__43055),
            .I(N__43049));
    LocalMux I__9585 (
            .O(N__43052),
            .I(N__43043));
    LocalMux I__9584 (
            .O(N__43049),
            .I(N__43043));
    InMux I__9583 (
            .O(N__43048),
            .I(N__43040));
    Span12Mux_v I__9582 (
            .O(N__43043),
            .I(N__43036));
    LocalMux I__9581 (
            .O(N__43040),
            .I(N__43033));
    InMux I__9580 (
            .O(N__43039),
            .I(N__43030));
    Odrv12 I__9579 (
            .O(N__43036),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv12 I__9578 (
            .O(N__43033),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__9577 (
            .O(N__43030),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__9576 (
            .O(N__43023),
            .I(N__43020));
    LocalMux I__9575 (
            .O(N__43020),
            .I(N__43017));
    Odrv12 I__9574 (
            .O(N__43017),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    CascadeMux I__9573 (
            .O(N__43014),
            .I(N__43010));
    CascadeMux I__9572 (
            .O(N__43013),
            .I(N__43007));
    InMux I__9571 (
            .O(N__43010),
            .I(N__43004));
    InMux I__9570 (
            .O(N__43007),
            .I(N__43001));
    LocalMux I__9569 (
            .O(N__43004),
            .I(N__42998));
    LocalMux I__9568 (
            .O(N__43001),
            .I(N__42994));
    Span4Mux_h I__9567 (
            .O(N__42998),
            .I(N__42991));
    InMux I__9566 (
            .O(N__42997),
            .I(N__42988));
    Span4Mux_h I__9565 (
            .O(N__42994),
            .I(N__42984));
    Span4Mux_v I__9564 (
            .O(N__42991),
            .I(N__42979));
    LocalMux I__9563 (
            .O(N__42988),
            .I(N__42979));
    InMux I__9562 (
            .O(N__42987),
            .I(N__42976));
    Odrv4 I__9561 (
            .O(N__42984),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__9560 (
            .O(N__42979),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__9559 (
            .O(N__42976),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__9558 (
            .O(N__42969),
            .I(N__42966));
    LocalMux I__9557 (
            .O(N__42966),
            .I(N__42963));
    Odrv4 I__9556 (
            .O(N__42963),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    CascadeMux I__9555 (
            .O(N__42960),
            .I(N__42956));
    CascadeMux I__9554 (
            .O(N__42959),
            .I(N__42953));
    InMux I__9553 (
            .O(N__42956),
            .I(N__42950));
    InMux I__9552 (
            .O(N__42953),
            .I(N__42947));
    LocalMux I__9551 (
            .O(N__42950),
            .I(N__42944));
    LocalMux I__9550 (
            .O(N__42947),
            .I(N__42941));
    Sp12to4 I__9549 (
            .O(N__42944),
            .I(N__42934));
    Span12Mux_h I__9548 (
            .O(N__42941),
            .I(N__42934));
    InMux I__9547 (
            .O(N__42940),
            .I(N__42931));
    InMux I__9546 (
            .O(N__42939),
            .I(N__42928));
    Odrv12 I__9545 (
            .O(N__42934),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__9544 (
            .O(N__42931),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__9543 (
            .O(N__42928),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__9542 (
            .O(N__42921),
            .I(N__42918));
    LocalMux I__9541 (
            .O(N__42918),
            .I(N__42915));
    Odrv4 I__9540 (
            .O(N__42915),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    CascadeMux I__9539 (
            .O(N__42912),
            .I(N__42909));
    InMux I__9538 (
            .O(N__42909),
            .I(N__42905));
    InMux I__9537 (
            .O(N__42908),
            .I(N__42902));
    LocalMux I__9536 (
            .O(N__42905),
            .I(N__42897));
    LocalMux I__9535 (
            .O(N__42902),
            .I(N__42897));
    Span4Mux_h I__9534 (
            .O(N__42897),
            .I(N__42892));
    InMux I__9533 (
            .O(N__42896),
            .I(N__42889));
    InMux I__9532 (
            .O(N__42895),
            .I(N__42886));
    Odrv4 I__9531 (
            .O(N__42892),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__9530 (
            .O(N__42889),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__9529 (
            .O(N__42886),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__9528 (
            .O(N__42879),
            .I(N__42876));
    LocalMux I__9527 (
            .O(N__42876),
            .I(N__42873));
    Odrv4 I__9526 (
            .O(N__42873),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    CascadeMux I__9525 (
            .O(N__42870),
            .I(N__42867));
    InMux I__9524 (
            .O(N__42867),
            .I(N__42863));
    InMux I__9523 (
            .O(N__42866),
            .I(N__42860));
    LocalMux I__9522 (
            .O(N__42863),
            .I(N__42856));
    LocalMux I__9521 (
            .O(N__42860),
            .I(N__42853));
    InMux I__9520 (
            .O(N__42859),
            .I(N__42850));
    Span4Mux_v I__9519 (
            .O(N__42856),
            .I(N__42845));
    Span4Mux_h I__9518 (
            .O(N__42853),
            .I(N__42845));
    LocalMux I__9517 (
            .O(N__42850),
            .I(N__42841));
    Span4Mux_v I__9516 (
            .O(N__42845),
            .I(N__42838));
    InMux I__9515 (
            .O(N__42844),
            .I(N__42835));
    Odrv12 I__9514 (
            .O(N__42841),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__9513 (
            .O(N__42838),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__9512 (
            .O(N__42835),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__9511 (
            .O(N__42828),
            .I(N__42825));
    LocalMux I__9510 (
            .O(N__42825),
            .I(N__42822));
    Odrv12 I__9509 (
            .O(N__42822),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__9508 (
            .O(N__42819),
            .I(N__42814));
    CascadeMux I__9507 (
            .O(N__42818),
            .I(N__42811));
    CascadeMux I__9506 (
            .O(N__42817),
            .I(N__42808));
    LocalMux I__9505 (
            .O(N__42814),
            .I(N__42805));
    InMux I__9504 (
            .O(N__42811),
            .I(N__42800));
    InMux I__9503 (
            .O(N__42808),
            .I(N__42800));
    Span4Mux_h I__9502 (
            .O(N__42805),
            .I(N__42794));
    LocalMux I__9501 (
            .O(N__42800),
            .I(N__42794));
    InMux I__9500 (
            .O(N__42799),
            .I(N__42791));
    Odrv4 I__9499 (
            .O(N__42794),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__9498 (
            .O(N__42791),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__9497 (
            .O(N__42786),
            .I(N__42783));
    LocalMux I__9496 (
            .O(N__42783),
            .I(N__42780));
    Odrv12 I__9495 (
            .O(N__42780),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__9494 (
            .O(N__42777),
            .I(N__42774));
    LocalMux I__9493 (
            .O(N__42774),
            .I(N__42771));
    Odrv4 I__9492 (
            .O(N__42771),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__9491 (
            .O(N__42768),
            .I(N__42765));
    LocalMux I__9490 (
            .O(N__42765),
            .I(N__42762));
    Odrv4 I__9489 (
            .O(N__42762),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__9488 (
            .O(N__42759),
            .I(N__42754));
    InMux I__9487 (
            .O(N__42758),
            .I(N__42751));
    CascadeMux I__9486 (
            .O(N__42757),
            .I(N__42748));
    LocalMux I__9485 (
            .O(N__42754),
            .I(N__42745));
    LocalMux I__9484 (
            .O(N__42751),
            .I(N__42742));
    InMux I__9483 (
            .O(N__42748),
            .I(N__42739));
    Sp12to4 I__9482 (
            .O(N__42745),
            .I(N__42731));
    Sp12to4 I__9481 (
            .O(N__42742),
            .I(N__42731));
    LocalMux I__9480 (
            .O(N__42739),
            .I(N__42731));
    InMux I__9479 (
            .O(N__42738),
            .I(N__42728));
    Odrv12 I__9478 (
            .O(N__42731),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__9477 (
            .O(N__42728),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__9476 (
            .O(N__42723),
            .I(N__42720));
    LocalMux I__9475 (
            .O(N__42720),
            .I(N__42717));
    Odrv12 I__9474 (
            .O(N__42717),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    CascadeMux I__9473 (
            .O(N__42714),
            .I(N__42710));
    CascadeMux I__9472 (
            .O(N__42713),
            .I(N__42707));
    InMux I__9471 (
            .O(N__42710),
            .I(N__42704));
    InMux I__9470 (
            .O(N__42707),
            .I(N__42701));
    LocalMux I__9469 (
            .O(N__42704),
            .I(N__42698));
    LocalMux I__9468 (
            .O(N__42701),
            .I(N__42694));
    Span4Mux_h I__9467 (
            .O(N__42698),
            .I(N__42691));
    InMux I__9466 (
            .O(N__42697),
            .I(N__42688));
    Span4Mux_v I__9465 (
            .O(N__42694),
            .I(N__42684));
    Sp12to4 I__9464 (
            .O(N__42691),
            .I(N__42679));
    LocalMux I__9463 (
            .O(N__42688),
            .I(N__42679));
    InMux I__9462 (
            .O(N__42687),
            .I(N__42676));
    Odrv4 I__9461 (
            .O(N__42684),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv12 I__9460 (
            .O(N__42679),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__9459 (
            .O(N__42676),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__9458 (
            .O(N__42669),
            .I(N__42666));
    LocalMux I__9457 (
            .O(N__42666),
            .I(N__42663));
    Span4Mux_v I__9456 (
            .O(N__42663),
            .I(N__42660));
    Odrv4 I__9455 (
            .O(N__42660),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__9454 (
            .O(N__42657),
            .I(N__42653));
    InMux I__9453 (
            .O(N__42656),
            .I(N__42650));
    LocalMux I__9452 (
            .O(N__42653),
            .I(N__42647));
    LocalMux I__9451 (
            .O(N__42650),
            .I(N__42644));
    Span4Mux_v I__9450 (
            .O(N__42647),
            .I(N__42641));
    Span4Mux_v I__9449 (
            .O(N__42644),
            .I(N__42637));
    Span4Mux_h I__9448 (
            .O(N__42641),
            .I(N__42634));
    InMux I__9447 (
            .O(N__42640),
            .I(N__42631));
    Span4Mux_v I__9446 (
            .O(N__42637),
            .I(N__42628));
    Odrv4 I__9445 (
            .O(N__42634),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9444 (
            .O(N__42631),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__9443 (
            .O(N__42628),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__9442 (
            .O(N__42621),
            .I(N__42618));
    LocalMux I__9441 (
            .O(N__42618),
            .I(N__42615));
    Odrv12 I__9440 (
            .O(N__42615),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    CascadeMux I__9439 (
            .O(N__42612),
            .I(N__42609));
    InMux I__9438 (
            .O(N__42609),
            .I(N__42606));
    LocalMux I__9437 (
            .O(N__42606),
            .I(N__42602));
    InMux I__9436 (
            .O(N__42605),
            .I(N__42599));
    Span4Mux_h I__9435 (
            .O(N__42602),
            .I(N__42593));
    LocalMux I__9434 (
            .O(N__42599),
            .I(N__42593));
    InMux I__9433 (
            .O(N__42598),
            .I(N__42590));
    Sp12to4 I__9432 (
            .O(N__42593),
            .I(N__42586));
    LocalMux I__9431 (
            .O(N__42590),
            .I(N__42583));
    InMux I__9430 (
            .O(N__42589),
            .I(N__42580));
    Odrv12 I__9429 (
            .O(N__42586),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__9428 (
            .O(N__42583),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__9427 (
            .O(N__42580),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__9426 (
            .O(N__42573),
            .I(N__42570));
    LocalMux I__9425 (
            .O(N__42570),
            .I(N__42567));
    Odrv4 I__9424 (
            .O(N__42567),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__9423 (
            .O(N__42564),
            .I(N__42561));
    LocalMux I__9422 (
            .O(N__42561),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__9421 (
            .O(N__42558),
            .I(N__42555));
    LocalMux I__9420 (
            .O(N__42555),
            .I(N__42552));
    Span4Mux_h I__9419 (
            .O(N__42552),
            .I(N__42547));
    InMux I__9418 (
            .O(N__42551),
            .I(N__42544));
    InMux I__9417 (
            .O(N__42550),
            .I(N__42541));
    Odrv4 I__9416 (
            .O(N__42547),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__9415 (
            .O(N__42544),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__9414 (
            .O(N__42541),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__9413 (
            .O(N__42534),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__9412 (
            .O(N__42531),
            .I(N__42528));
    LocalMux I__9411 (
            .O(N__42528),
            .I(N__42525));
    Span4Mux_h I__9410 (
            .O(N__42525),
            .I(N__42522));
    Odrv4 I__9409 (
            .O(N__42522),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__9408 (
            .O(N__42519),
            .I(N__42516));
    LocalMux I__9407 (
            .O(N__42516),
            .I(N__42512));
    InMux I__9406 (
            .O(N__42515),
            .I(N__42509));
    Span4Mux_v I__9405 (
            .O(N__42512),
            .I(N__42505));
    LocalMux I__9404 (
            .O(N__42509),
            .I(N__42502));
    InMux I__9403 (
            .O(N__42508),
            .I(N__42499));
    Odrv4 I__9402 (
            .O(N__42505),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__9401 (
            .O(N__42502),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__9400 (
            .O(N__42499),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__9399 (
            .O(N__42492),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__9398 (
            .O(N__42489),
            .I(N__42486));
    LocalMux I__9397 (
            .O(N__42486),
            .I(N__42482));
    InMux I__9396 (
            .O(N__42485),
            .I(N__42479));
    Span4Mux_v I__9395 (
            .O(N__42482),
            .I(N__42473));
    LocalMux I__9394 (
            .O(N__42479),
            .I(N__42473));
    InMux I__9393 (
            .O(N__42478),
            .I(N__42470));
    Odrv4 I__9392 (
            .O(N__42473),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__9391 (
            .O(N__42470),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__9390 (
            .O(N__42465),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__9389 (
            .O(N__42462),
            .I(bfn_17_18_0_));
    InMux I__9388 (
            .O(N__42459),
            .I(N__42454));
    InMux I__9387 (
            .O(N__42458),
            .I(N__42451));
    InMux I__9386 (
            .O(N__42457),
            .I(N__42448));
    LocalMux I__9385 (
            .O(N__42454),
            .I(N__42445));
    LocalMux I__9384 (
            .O(N__42451),
            .I(N__42442));
    LocalMux I__9383 (
            .O(N__42448),
            .I(N__42439));
    Span4Mux_h I__9382 (
            .O(N__42445),
            .I(N__42436));
    Span4Mux_v I__9381 (
            .O(N__42442),
            .I(N__42431));
    Span4Mux_h I__9380 (
            .O(N__42439),
            .I(N__42431));
    Span4Mux_v I__9379 (
            .O(N__42436),
            .I(N__42428));
    Odrv4 I__9378 (
            .O(N__42431),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__9377 (
            .O(N__42428),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__9376 (
            .O(N__42423),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__9375 (
            .O(N__42420),
            .I(N__42415));
    InMux I__9374 (
            .O(N__42419),
            .I(N__42412));
    InMux I__9373 (
            .O(N__42418),
            .I(N__42409));
    LocalMux I__9372 (
            .O(N__42415),
            .I(N__42406));
    LocalMux I__9371 (
            .O(N__42412),
            .I(N__42401));
    LocalMux I__9370 (
            .O(N__42409),
            .I(N__42401));
    Span4Mux_v I__9369 (
            .O(N__42406),
            .I(N__42398));
    Odrv4 I__9368 (
            .O(N__42401),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__9367 (
            .O(N__42398),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__9366 (
            .O(N__42393),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__9365 (
            .O(N__42390),
            .I(N__42385));
    InMux I__9364 (
            .O(N__42389),
            .I(N__42382));
    InMux I__9363 (
            .O(N__42388),
            .I(N__42379));
    LocalMux I__9362 (
            .O(N__42385),
            .I(N__42376));
    LocalMux I__9361 (
            .O(N__42382),
            .I(N__42373));
    LocalMux I__9360 (
            .O(N__42379),
            .I(N__42370));
    Span4Mux_h I__9359 (
            .O(N__42376),
            .I(N__42367));
    Span4Mux_h I__9358 (
            .O(N__42373),
            .I(N__42362));
    Span4Mux_v I__9357 (
            .O(N__42370),
            .I(N__42362));
    Odrv4 I__9356 (
            .O(N__42367),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__9355 (
            .O(N__42362),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__9354 (
            .O(N__42357),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__9353 (
            .O(N__42354),
            .I(N__42349));
    InMux I__9352 (
            .O(N__42353),
            .I(N__42346));
    InMux I__9351 (
            .O(N__42352),
            .I(N__42343));
    LocalMux I__9350 (
            .O(N__42349),
            .I(N__42340));
    LocalMux I__9349 (
            .O(N__42346),
            .I(N__42337));
    LocalMux I__9348 (
            .O(N__42343),
            .I(N__42334));
    Span4Mux_v I__9347 (
            .O(N__42340),
            .I(N__42331));
    Odrv4 I__9346 (
            .O(N__42337),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__9345 (
            .O(N__42334),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__9344 (
            .O(N__42331),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__9343 (
            .O(N__42324),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__9342 (
            .O(N__42321),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__9341 (
            .O(N__42318),
            .I(N__42315));
    InMux I__9340 (
            .O(N__42315),
            .I(N__42311));
    InMux I__9339 (
            .O(N__42314),
            .I(N__42307));
    LocalMux I__9338 (
            .O(N__42311),
            .I(N__42304));
    InMux I__9337 (
            .O(N__42310),
            .I(N__42301));
    LocalMux I__9336 (
            .O(N__42307),
            .I(N__42298));
    Span4Mux_h I__9335 (
            .O(N__42304),
            .I(N__42295));
    LocalMux I__9334 (
            .O(N__42301),
            .I(N__42292));
    Sp12to4 I__9333 (
            .O(N__42298),
            .I(N__42289));
    Odrv4 I__9332 (
            .O(N__42295),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv4 I__9331 (
            .O(N__42292),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv12 I__9330 (
            .O(N__42289),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    InMux I__9329 (
            .O(N__42282),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__9328 (
            .O(N__42279),
            .I(N__42275));
    CascadeMux I__9327 (
            .O(N__42278),
            .I(N__42272));
    LocalMux I__9326 (
            .O(N__42275),
            .I(N__42269));
    InMux I__9325 (
            .O(N__42272),
            .I(N__42265));
    Span4Mux_h I__9324 (
            .O(N__42269),
            .I(N__42262));
    InMux I__9323 (
            .O(N__42268),
            .I(N__42259));
    LocalMux I__9322 (
            .O(N__42265),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__9321 (
            .O(N__42262),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__9320 (
            .O(N__42259),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__9319 (
            .O(N__42252),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__9318 (
            .O(N__42249),
            .I(N__42245));
    CascadeMux I__9317 (
            .O(N__42248),
            .I(N__42242));
    LocalMux I__9316 (
            .O(N__42245),
            .I(N__42239));
    InMux I__9315 (
            .O(N__42242),
            .I(N__42236));
    Span4Mux_v I__9314 (
            .O(N__42239),
            .I(N__42230));
    LocalMux I__9313 (
            .O(N__42236),
            .I(N__42230));
    InMux I__9312 (
            .O(N__42235),
            .I(N__42227));
    Odrv4 I__9311 (
            .O(N__42230),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__9310 (
            .O(N__42227),
            .I(\current_shift_inst.un4_control_input1_17 ));
    InMux I__9309 (
            .O(N__42222),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__9308 (
            .O(N__42219),
            .I(N__42216));
    LocalMux I__9307 (
            .O(N__42216),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__9306 (
            .O(N__42213),
            .I(N__42208));
    InMux I__9305 (
            .O(N__42212),
            .I(N__42205));
    InMux I__9304 (
            .O(N__42211),
            .I(N__42202));
    LocalMux I__9303 (
            .O(N__42208),
            .I(N__42199));
    LocalMux I__9302 (
            .O(N__42205),
            .I(N__42196));
    LocalMux I__9301 (
            .O(N__42202),
            .I(N__42193));
    Span4Mux_h I__9300 (
            .O(N__42199),
            .I(N__42188));
    Span4Mux_v I__9299 (
            .O(N__42196),
            .I(N__42188));
    Odrv12 I__9298 (
            .O(N__42193),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__9297 (
            .O(N__42188),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__9296 (
            .O(N__42183),
            .I(bfn_17_17_0_));
    CascadeMux I__9295 (
            .O(N__42180),
            .I(N__42177));
    InMux I__9294 (
            .O(N__42177),
            .I(N__42172));
    InMux I__9293 (
            .O(N__42176),
            .I(N__42169));
    InMux I__9292 (
            .O(N__42175),
            .I(N__42166));
    LocalMux I__9291 (
            .O(N__42172),
            .I(N__42163));
    LocalMux I__9290 (
            .O(N__42169),
            .I(N__42160));
    LocalMux I__9289 (
            .O(N__42166),
            .I(N__42157));
    Span4Mux_h I__9288 (
            .O(N__42163),
            .I(N__42152));
    Span4Mux_v I__9287 (
            .O(N__42160),
            .I(N__42152));
    Span4Mux_v I__9286 (
            .O(N__42157),
            .I(N__42149));
    Odrv4 I__9285 (
            .O(N__42152),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__9284 (
            .O(N__42149),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__9283 (
            .O(N__42144),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    CascadeMux I__9282 (
            .O(N__42141),
            .I(N__42137));
    InMux I__9281 (
            .O(N__42140),
            .I(N__42133));
    InMux I__9280 (
            .O(N__42137),
            .I(N__42130));
    InMux I__9279 (
            .O(N__42136),
            .I(N__42127));
    LocalMux I__9278 (
            .O(N__42133),
            .I(N__42124));
    LocalMux I__9277 (
            .O(N__42130),
            .I(N__42121));
    LocalMux I__9276 (
            .O(N__42127),
            .I(N__42118));
    Span4Mux_h I__9275 (
            .O(N__42124),
            .I(N__42113));
    Span4Mux_v I__9274 (
            .O(N__42121),
            .I(N__42113));
    Span4Mux_v I__9273 (
            .O(N__42118),
            .I(N__42110));
    Odrv4 I__9272 (
            .O(N__42113),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__9271 (
            .O(N__42110),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__9270 (
            .O(N__42105),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__9269 (
            .O(N__42102),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__9268 (
            .O(N__42099),
            .I(N__42096));
    LocalMux I__9267 (
            .O(N__42096),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    CascadeMux I__9266 (
            .O(N__42093),
            .I(N__42090));
    InMux I__9265 (
            .O(N__42090),
            .I(N__42086));
    InMux I__9264 (
            .O(N__42089),
            .I(N__42082));
    LocalMux I__9263 (
            .O(N__42086),
            .I(N__42079));
    InMux I__9262 (
            .O(N__42085),
            .I(N__42076));
    LocalMux I__9261 (
            .O(N__42082),
            .I(N__42073));
    Span4Mux_h I__9260 (
            .O(N__42079),
            .I(N__42068));
    LocalMux I__9259 (
            .O(N__42076),
            .I(N__42068));
    Span4Mux_v I__9258 (
            .O(N__42073),
            .I(N__42065));
    Odrv4 I__9257 (
            .O(N__42068),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__9256 (
            .O(N__42065),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__9255 (
            .O(N__42060),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__9254 (
            .O(N__42057),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__9253 (
            .O(N__42054),
            .I(N__42050));
    InMux I__9252 (
            .O(N__42053),
            .I(N__42047));
    LocalMux I__9251 (
            .O(N__42050),
            .I(N__42044));
    LocalMux I__9250 (
            .O(N__42047),
            .I(N__42041));
    Span4Mux_v I__9249 (
            .O(N__42044),
            .I(N__42037));
    Span4Mux_h I__9248 (
            .O(N__42041),
            .I(N__42034));
    InMux I__9247 (
            .O(N__42040),
            .I(N__42031));
    Odrv4 I__9246 (
            .O(N__42037),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__9245 (
            .O(N__42034),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__9244 (
            .O(N__42031),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__9243 (
            .O(N__42024),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__9242 (
            .O(N__42021),
            .I(N__42018));
    LocalMux I__9241 (
            .O(N__42018),
            .I(N__42015));
    Span4Mux_h I__9240 (
            .O(N__42015),
            .I(N__42012));
    Odrv4 I__9239 (
            .O(N__42012),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__9238 (
            .O(N__42009),
            .I(N__42005));
    InMux I__9237 (
            .O(N__42008),
            .I(N__42002));
    LocalMux I__9236 (
            .O(N__42005),
            .I(N__41999));
    LocalMux I__9235 (
            .O(N__42002),
            .I(N__41996));
    Span4Mux_h I__9234 (
            .O(N__41999),
            .I(N__41992));
    Span4Mux_h I__9233 (
            .O(N__41996),
            .I(N__41989));
    InMux I__9232 (
            .O(N__41995),
            .I(N__41986));
    Odrv4 I__9231 (
            .O(N__41992),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__9230 (
            .O(N__41989),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__9229 (
            .O(N__41986),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__9228 (
            .O(N__41979),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__9227 (
            .O(N__41976),
            .I(N__41973));
    LocalMux I__9226 (
            .O(N__41973),
            .I(N__41969));
    InMux I__9225 (
            .O(N__41972),
            .I(N__41966));
    Span4Mux_v I__9224 (
            .O(N__41969),
            .I(N__41960));
    LocalMux I__9223 (
            .O(N__41966),
            .I(N__41960));
    InMux I__9222 (
            .O(N__41965),
            .I(N__41957));
    Odrv4 I__9221 (
            .O(N__41960),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__9220 (
            .O(N__41957),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__9219 (
            .O(N__41952),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__9218 (
            .O(N__41949),
            .I(N__41946));
    LocalMux I__9217 (
            .O(N__41946),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__9216 (
            .O(N__41943),
            .I(N__41940));
    LocalMux I__9215 (
            .O(N__41940),
            .I(N__41937));
    Span4Mux_v I__9214 (
            .O(N__41937),
            .I(N__41932));
    InMux I__9213 (
            .O(N__41936),
            .I(N__41929));
    InMux I__9212 (
            .O(N__41935),
            .I(N__41926));
    Odrv4 I__9211 (
            .O(N__41932),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__9210 (
            .O(N__41929),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__9209 (
            .O(N__41926),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__9208 (
            .O(N__41919),
            .I(bfn_17_16_0_));
    InMux I__9207 (
            .O(N__41916),
            .I(N__41913));
    LocalMux I__9206 (
            .O(N__41913),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__9205 (
            .O(N__41910),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__9204 (
            .O(N__41907),
            .I(N__41904));
    LocalMux I__9203 (
            .O(N__41904),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__9202 (
            .O(N__41901),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__9201 (
            .O(N__41898),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__9200 (
            .O(N__41895),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__9199 (
            .O(N__41892),
            .I(N__41889));
    LocalMux I__9198 (
            .O(N__41889),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__9197 (
            .O(N__41886),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    CascadeMux I__9196 (
            .O(N__41883),
            .I(N__41879));
    InMux I__9195 (
            .O(N__41882),
            .I(N__41876));
    InMux I__9194 (
            .O(N__41879),
            .I(N__41873));
    LocalMux I__9193 (
            .O(N__41876),
            .I(N__41870));
    LocalMux I__9192 (
            .O(N__41873),
            .I(N__41867));
    Span4Mux_h I__9191 (
            .O(N__41870),
            .I(N__41864));
    Span4Mux_h I__9190 (
            .O(N__41867),
            .I(N__41861));
    Span4Mux_v I__9189 (
            .O(N__41864),
            .I(N__41856));
    Span4Mux_h I__9188 (
            .O(N__41861),
            .I(N__41856));
    Odrv4 I__9187 (
            .O(N__41856),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__9186 (
            .O(N__41853),
            .I(N__41850));
    InMux I__9185 (
            .O(N__41850),
            .I(N__41847));
    LocalMux I__9184 (
            .O(N__41847),
            .I(N__41844));
    Span4Mux_h I__9183 (
            .O(N__41844),
            .I(N__41841));
    Odrv4 I__9182 (
            .O(N__41841),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__9181 (
            .O(N__41838),
            .I(N__41833));
    InMux I__9180 (
            .O(N__41837),
            .I(N__41828));
    InMux I__9179 (
            .O(N__41836),
            .I(N__41828));
    LocalMux I__9178 (
            .O(N__41833),
            .I(N__41824));
    LocalMux I__9177 (
            .O(N__41828),
            .I(N__41821));
    InMux I__9176 (
            .O(N__41827),
            .I(N__41818));
    Span4Mux_v I__9175 (
            .O(N__41824),
            .I(N__41815));
    Span4Mux_v I__9174 (
            .O(N__41821),
            .I(N__41812));
    LocalMux I__9173 (
            .O(N__41818),
            .I(N__41809));
    Odrv4 I__9172 (
            .O(N__41815),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__9171 (
            .O(N__41812),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__9170 (
            .O(N__41809),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    CascadeMux I__9169 (
            .O(N__41802),
            .I(N__41799));
    InMux I__9168 (
            .O(N__41799),
            .I(N__41796));
    LocalMux I__9167 (
            .O(N__41796),
            .I(N__41793));
    Span4Mux_h I__9166 (
            .O(N__41793),
            .I(N__41790));
    Odrv4 I__9165 (
            .O(N__41790),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ));
    InMux I__9164 (
            .O(N__41787),
            .I(N__41784));
    LocalMux I__9163 (
            .O(N__41784),
            .I(N__41781));
    Odrv4 I__9162 (
            .O(N__41781),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__9161 (
            .O(N__41778),
            .I(N__41775));
    LocalMux I__9160 (
            .O(N__41775),
            .I(N__41771));
    InMux I__9159 (
            .O(N__41774),
            .I(N__41768));
    Span4Mux_v I__9158 (
            .O(N__41771),
            .I(N__41762));
    LocalMux I__9157 (
            .O(N__41768),
            .I(N__41762));
    InMux I__9156 (
            .O(N__41767),
            .I(N__41759));
    Odrv4 I__9155 (
            .O(N__41762),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__9154 (
            .O(N__41759),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__9153 (
            .O(N__41754),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__9152 (
            .O(N__41751),
            .I(N__41748));
    LocalMux I__9151 (
            .O(N__41748),
            .I(N__41745));
    Span4Mux_v I__9150 (
            .O(N__41745),
            .I(N__41740));
    InMux I__9149 (
            .O(N__41744),
            .I(N__41737));
    InMux I__9148 (
            .O(N__41743),
            .I(N__41734));
    Odrv4 I__9147 (
            .O(N__41740),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__9146 (
            .O(N__41737),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__9145 (
            .O(N__41734),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__9144 (
            .O(N__41727),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__9143 (
            .O(N__41724),
            .I(N__41721));
    LocalMux I__9142 (
            .O(N__41721),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__9141 (
            .O(N__41718),
            .I(N__41713));
    InMux I__9140 (
            .O(N__41717),
            .I(N__41708));
    InMux I__9139 (
            .O(N__41716),
            .I(N__41708));
    LocalMux I__9138 (
            .O(N__41713),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__9137 (
            .O(N__41708),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__9136 (
            .O(N__41703),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    CascadeMux I__9135 (
            .O(N__41700),
            .I(N__41697));
    InMux I__9134 (
            .O(N__41697),
            .I(N__41692));
    InMux I__9133 (
            .O(N__41696),
            .I(N__41687));
    InMux I__9132 (
            .O(N__41695),
            .I(N__41687));
    LocalMux I__9131 (
            .O(N__41692),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__9130 (
            .O(N__41687),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__9129 (
            .O(N__41682),
            .I(N__41679));
    LocalMux I__9128 (
            .O(N__41679),
            .I(N__41673));
    InMux I__9127 (
            .O(N__41678),
            .I(N__41670));
    InMux I__9126 (
            .O(N__41677),
            .I(N__41665));
    InMux I__9125 (
            .O(N__41676),
            .I(N__41665));
    Span4Mux_h I__9124 (
            .O(N__41673),
            .I(N__41662));
    LocalMux I__9123 (
            .O(N__41670),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__9122 (
            .O(N__41665),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    Odrv4 I__9121 (
            .O(N__41662),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__9120 (
            .O(N__41655),
            .I(N__41652));
    LocalMux I__9119 (
            .O(N__41652),
            .I(N__41648));
    InMux I__9118 (
            .O(N__41651),
            .I(N__41645));
    Odrv4 I__9117 (
            .O(N__41648),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    LocalMux I__9116 (
            .O(N__41645),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__9115 (
            .O(N__41640),
            .I(N__41634));
    InMux I__9114 (
            .O(N__41639),
            .I(N__41634));
    LocalMux I__9113 (
            .O(N__41634),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    InMux I__9112 (
            .O(N__41631),
            .I(N__41625));
    InMux I__9111 (
            .O(N__41630),
            .I(N__41625));
    LocalMux I__9110 (
            .O(N__41625),
            .I(N__41620));
    InMux I__9109 (
            .O(N__41624),
            .I(N__41617));
    InMux I__9108 (
            .O(N__41623),
            .I(N__41614));
    Span4Mux_v I__9107 (
            .O(N__41620),
            .I(N__41609));
    LocalMux I__9106 (
            .O(N__41617),
            .I(N__41609));
    LocalMux I__9105 (
            .O(N__41614),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__9104 (
            .O(N__41609),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__9103 (
            .O(N__41604),
            .I(N__41601));
    LocalMux I__9102 (
            .O(N__41601),
            .I(N__41598));
    Span4Mux_h I__9101 (
            .O(N__41598),
            .I(N__41594));
    InMux I__9100 (
            .O(N__41597),
            .I(N__41591));
    Odrv4 I__9099 (
            .O(N__41594),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    LocalMux I__9098 (
            .O(N__41591),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__9097 (
            .O(N__41586),
            .I(N__41582));
    InMux I__9096 (
            .O(N__41585),
            .I(N__41579));
    LocalMux I__9095 (
            .O(N__41582),
            .I(N__41576));
    LocalMux I__9094 (
            .O(N__41579),
            .I(N__41570));
    Sp12to4 I__9093 (
            .O(N__41576),
            .I(N__41570));
    InMux I__9092 (
            .O(N__41575),
            .I(N__41567));
    Span12Mux_s10_h I__9091 (
            .O(N__41570),
            .I(N__41564));
    LocalMux I__9090 (
            .O(N__41567),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    Odrv12 I__9089 (
            .O(N__41564),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    InMux I__9088 (
            .O(N__41559),
            .I(N__41555));
    InMux I__9087 (
            .O(N__41558),
            .I(N__41552));
    LocalMux I__9086 (
            .O(N__41555),
            .I(N__41547));
    LocalMux I__9085 (
            .O(N__41552),
            .I(N__41544));
    InMux I__9084 (
            .O(N__41551),
            .I(N__41541));
    InMux I__9083 (
            .O(N__41550),
            .I(N__41538));
    Span4Mux_v I__9082 (
            .O(N__41547),
            .I(N__41533));
    Span4Mux_h I__9081 (
            .O(N__41544),
            .I(N__41533));
    LocalMux I__9080 (
            .O(N__41541),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__9079 (
            .O(N__41538),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv4 I__9078 (
            .O(N__41533),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__9077 (
            .O(N__41526),
            .I(N__41522));
    InMux I__9076 (
            .O(N__41525),
            .I(N__41519));
    LocalMux I__9075 (
            .O(N__41522),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    LocalMux I__9074 (
            .O(N__41519),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    InMux I__9073 (
            .O(N__41514),
            .I(N__41510));
    InMux I__9072 (
            .O(N__41513),
            .I(N__41506));
    LocalMux I__9071 (
            .O(N__41510),
            .I(N__41503));
    InMux I__9070 (
            .O(N__41509),
            .I(N__41500));
    LocalMux I__9069 (
            .O(N__41506),
            .I(N__41497));
    Span4Mux_v I__9068 (
            .O(N__41503),
            .I(N__41493));
    LocalMux I__9067 (
            .O(N__41500),
            .I(N__41490));
    Span4Mux_v I__9066 (
            .O(N__41497),
            .I(N__41487));
    InMux I__9065 (
            .O(N__41496),
            .I(N__41484));
    Odrv4 I__9064 (
            .O(N__41493),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    Odrv4 I__9063 (
            .O(N__41490),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    Odrv4 I__9062 (
            .O(N__41487),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__9061 (
            .O(N__41484),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__9060 (
            .O(N__41475),
            .I(N__41471));
    InMux I__9059 (
            .O(N__41474),
            .I(N__41468));
    LocalMux I__9058 (
            .O(N__41471),
            .I(N__41465));
    LocalMux I__9057 (
            .O(N__41468),
            .I(N__41462));
    Span4Mux_h I__9056 (
            .O(N__41465),
            .I(N__41456));
    Span4Mux_v I__9055 (
            .O(N__41462),
            .I(N__41456));
    InMux I__9054 (
            .O(N__41461),
            .I(N__41453));
    Span4Mux_v I__9053 (
            .O(N__41456),
            .I(N__41450));
    LocalMux I__9052 (
            .O(N__41453),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv4 I__9051 (
            .O(N__41450),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    CascadeMux I__9050 (
            .O(N__41445),
            .I(N__41442));
    InMux I__9049 (
            .O(N__41442),
            .I(N__41439));
    LocalMux I__9048 (
            .O(N__41439),
            .I(N__41436));
    Odrv12 I__9047 (
            .O(N__41436),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    InMux I__9046 (
            .O(N__41433),
            .I(N__41427));
    InMux I__9045 (
            .O(N__41432),
            .I(N__41424));
    InMux I__9044 (
            .O(N__41431),
            .I(N__41421));
    InMux I__9043 (
            .O(N__41430),
            .I(N__41418));
    LocalMux I__9042 (
            .O(N__41427),
            .I(N__41413));
    LocalMux I__9041 (
            .O(N__41424),
            .I(N__41413));
    LocalMux I__9040 (
            .O(N__41421),
            .I(N__41408));
    LocalMux I__9039 (
            .O(N__41418),
            .I(N__41408));
    Span4Mux_v I__9038 (
            .O(N__41413),
            .I(N__41405));
    Odrv4 I__9037 (
            .O(N__41408),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__9036 (
            .O(N__41405),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__9035 (
            .O(N__41400),
            .I(N__41397));
    LocalMux I__9034 (
            .O(N__41397),
            .I(N__41392));
    InMux I__9033 (
            .O(N__41396),
            .I(N__41389));
    InMux I__9032 (
            .O(N__41395),
            .I(N__41386));
    Span4Mux_h I__9031 (
            .O(N__41392),
            .I(N__41383));
    LocalMux I__9030 (
            .O(N__41389),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    LocalMux I__9029 (
            .O(N__41386),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv4 I__9028 (
            .O(N__41383),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    InMux I__9027 (
            .O(N__41376),
            .I(N__41371));
    InMux I__9026 (
            .O(N__41375),
            .I(N__41368));
    InMux I__9025 (
            .O(N__41374),
            .I(N__41364));
    LocalMux I__9024 (
            .O(N__41371),
            .I(N__41359));
    LocalMux I__9023 (
            .O(N__41368),
            .I(N__41359));
    InMux I__9022 (
            .O(N__41367),
            .I(N__41356));
    LocalMux I__9021 (
            .O(N__41364),
            .I(N__41353));
    Span4Mux_v I__9020 (
            .O(N__41359),
            .I(N__41350));
    LocalMux I__9019 (
            .O(N__41356),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__9018 (
            .O(N__41353),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__9017 (
            .O(N__41350),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__9016 (
            .O(N__41343),
            .I(N__41338));
    InMux I__9015 (
            .O(N__41342),
            .I(N__41335));
    InMux I__9014 (
            .O(N__41341),
            .I(N__41332));
    LocalMux I__9013 (
            .O(N__41338),
            .I(N__41329));
    LocalMux I__9012 (
            .O(N__41335),
            .I(N__41326));
    LocalMux I__9011 (
            .O(N__41332),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv12 I__9010 (
            .O(N__41329),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv4 I__9009 (
            .O(N__41326),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    CascadeMux I__9008 (
            .O(N__41319),
            .I(N__41315));
    InMux I__9007 (
            .O(N__41318),
            .I(N__41312));
    InMux I__9006 (
            .O(N__41315),
            .I(N__41309));
    LocalMux I__9005 (
            .O(N__41312),
            .I(N__41305));
    LocalMux I__9004 (
            .O(N__41309),
            .I(N__41302));
    InMux I__9003 (
            .O(N__41308),
            .I(N__41299));
    Span4Mux_v I__9002 (
            .O(N__41305),
            .I(N__41294));
    Span4Mux_h I__9001 (
            .O(N__41302),
            .I(N__41294));
    LocalMux I__9000 (
            .O(N__41299),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__8999 (
            .O(N__41294),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__8998 (
            .O(N__41289),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    IoInMux I__8997 (
            .O(N__41286),
            .I(N__41283));
    LocalMux I__8996 (
            .O(N__41283),
            .I(N__41280));
    IoSpan4Mux I__8995 (
            .O(N__41280),
            .I(N__41266));
    InMux I__8994 (
            .O(N__41279),
            .I(N__41254));
    InMux I__8993 (
            .O(N__41278),
            .I(N__41254));
    InMux I__8992 (
            .O(N__41277),
            .I(N__41254));
    InMux I__8991 (
            .O(N__41276),
            .I(N__41254));
    InMux I__8990 (
            .O(N__41275),
            .I(N__41235));
    InMux I__8989 (
            .O(N__41274),
            .I(N__41235));
    InMux I__8988 (
            .O(N__41273),
            .I(N__41235));
    InMux I__8987 (
            .O(N__41272),
            .I(N__41226));
    InMux I__8986 (
            .O(N__41271),
            .I(N__41226));
    InMux I__8985 (
            .O(N__41270),
            .I(N__41226));
    InMux I__8984 (
            .O(N__41269),
            .I(N__41226));
    Sp12to4 I__8983 (
            .O(N__41266),
            .I(N__41223));
    InMux I__8982 (
            .O(N__41265),
            .I(N__41216));
    InMux I__8981 (
            .O(N__41264),
            .I(N__41216));
    InMux I__8980 (
            .O(N__41263),
            .I(N__41216));
    LocalMux I__8979 (
            .O(N__41254),
            .I(N__41208));
    InMux I__8978 (
            .O(N__41253),
            .I(N__41199));
    InMux I__8977 (
            .O(N__41252),
            .I(N__41199));
    InMux I__8976 (
            .O(N__41251),
            .I(N__41199));
    InMux I__8975 (
            .O(N__41250),
            .I(N__41199));
    InMux I__8974 (
            .O(N__41249),
            .I(N__41190));
    InMux I__8973 (
            .O(N__41248),
            .I(N__41190));
    InMux I__8972 (
            .O(N__41247),
            .I(N__41190));
    InMux I__8971 (
            .O(N__41246),
            .I(N__41190));
    InMux I__8970 (
            .O(N__41245),
            .I(N__41181));
    InMux I__8969 (
            .O(N__41244),
            .I(N__41181));
    InMux I__8968 (
            .O(N__41243),
            .I(N__41181));
    InMux I__8967 (
            .O(N__41242),
            .I(N__41181));
    LocalMux I__8966 (
            .O(N__41235),
            .I(N__41178));
    LocalMux I__8965 (
            .O(N__41226),
            .I(N__41175));
    Span12Mux_v I__8964 (
            .O(N__41223),
            .I(N__41172));
    LocalMux I__8963 (
            .O(N__41216),
            .I(N__41169));
    InMux I__8962 (
            .O(N__41215),
            .I(N__41166));
    InMux I__8961 (
            .O(N__41214),
            .I(N__41157));
    InMux I__8960 (
            .O(N__41213),
            .I(N__41157));
    InMux I__8959 (
            .O(N__41212),
            .I(N__41157));
    InMux I__8958 (
            .O(N__41211),
            .I(N__41157));
    Span4Mux_h I__8957 (
            .O(N__41208),
            .I(N__41144));
    LocalMux I__8956 (
            .O(N__41199),
            .I(N__41144));
    LocalMux I__8955 (
            .O(N__41190),
            .I(N__41144));
    LocalMux I__8954 (
            .O(N__41181),
            .I(N__41144));
    Span4Mux_v I__8953 (
            .O(N__41178),
            .I(N__41144));
    Span4Mux_v I__8952 (
            .O(N__41175),
            .I(N__41144));
    Span12Mux_v I__8951 (
            .O(N__41172),
            .I(N__41141));
    Odrv4 I__8950 (
            .O(N__41169),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__8949 (
            .O(N__41166),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__8948 (
            .O(N__41157),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__8947 (
            .O(N__41144),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__8946 (
            .O(N__41141),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__8945 (
            .O(N__41130),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__8944 (
            .O(N__41127),
            .I(N__41124));
    InMux I__8943 (
            .O(N__41124),
            .I(N__41121));
    LocalMux I__8942 (
            .O(N__41121),
            .I(N__41116));
    InMux I__8941 (
            .O(N__41120),
            .I(N__41113));
    InMux I__8940 (
            .O(N__41119),
            .I(N__41110));
    Span4Mux_h I__8939 (
            .O(N__41116),
            .I(N__41107));
    LocalMux I__8938 (
            .O(N__41113),
            .I(N__41104));
    LocalMux I__8937 (
            .O(N__41110),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__8936 (
            .O(N__41107),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv12 I__8935 (
            .O(N__41104),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__8934 (
            .O(N__41097),
            .I(N__41094));
    InMux I__8933 (
            .O(N__41094),
            .I(N__41091));
    LocalMux I__8932 (
            .O(N__41091),
            .I(N__41088));
    Span4Mux_h I__8931 (
            .O(N__41088),
            .I(N__41085));
    Odrv4 I__8930 (
            .O(N__41085),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    CascadeMux I__8929 (
            .O(N__41082),
            .I(N__41078));
    InMux I__8928 (
            .O(N__41081),
            .I(N__41072));
    InMux I__8927 (
            .O(N__41078),
            .I(N__41072));
    InMux I__8926 (
            .O(N__41077),
            .I(N__41069));
    LocalMux I__8925 (
            .O(N__41072),
            .I(N__41066));
    LocalMux I__8924 (
            .O(N__41069),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__8923 (
            .O(N__41066),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    CascadeMux I__8922 (
            .O(N__41061),
            .I(N__41058));
    InMux I__8921 (
            .O(N__41058),
            .I(N__41053));
    InMux I__8920 (
            .O(N__41057),
            .I(N__41050));
    InMux I__8919 (
            .O(N__41056),
            .I(N__41047));
    LocalMux I__8918 (
            .O(N__41053),
            .I(N__41042));
    LocalMux I__8917 (
            .O(N__41050),
            .I(N__41042));
    LocalMux I__8916 (
            .O(N__41047),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__8915 (
            .O(N__41042),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__8914 (
            .O(N__41037),
            .I(N__41034));
    LocalMux I__8913 (
            .O(N__41034),
            .I(N__41031));
    Odrv4 I__8912 (
            .O(N__41031),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    InMux I__8911 (
            .O(N__41028),
            .I(N__41025));
    LocalMux I__8910 (
            .O(N__41025),
            .I(N__41020));
    InMux I__8909 (
            .O(N__41024),
            .I(N__41017));
    InMux I__8908 (
            .O(N__41023),
            .I(N__41014));
    Span4Mux_h I__8907 (
            .O(N__41020),
            .I(N__41011));
    LocalMux I__8906 (
            .O(N__41017),
            .I(N__41008));
    LocalMux I__8905 (
            .O(N__41014),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    Odrv4 I__8904 (
            .O(N__41011),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    Odrv4 I__8903 (
            .O(N__41008),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    InMux I__8902 (
            .O(N__41001),
            .I(N__40998));
    LocalMux I__8901 (
            .O(N__40998),
            .I(N__40993));
    InMux I__8900 (
            .O(N__40997),
            .I(N__40988));
    InMux I__8899 (
            .O(N__40996),
            .I(N__40988));
    Span4Mux_h I__8898 (
            .O(N__40993),
            .I(N__40982));
    LocalMux I__8897 (
            .O(N__40988),
            .I(N__40982));
    InMux I__8896 (
            .O(N__40987),
            .I(N__40979));
    Span4Mux_v I__8895 (
            .O(N__40982),
            .I(N__40976));
    LocalMux I__8894 (
            .O(N__40979),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    Odrv4 I__8893 (
            .O(N__40976),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__8892 (
            .O(N__40971),
            .I(N__40968));
    LocalMux I__8891 (
            .O(N__40968),
            .I(N__40965));
    Odrv4 I__8890 (
            .O(N__40965),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__8889 (
            .O(N__40962),
            .I(N__40957));
    InMux I__8888 (
            .O(N__40961),
            .I(N__40954));
    InMux I__8887 (
            .O(N__40960),
            .I(N__40951));
    InMux I__8886 (
            .O(N__40957),
            .I(N__40948));
    LocalMux I__8885 (
            .O(N__40954),
            .I(N__40940));
    LocalMux I__8884 (
            .O(N__40951),
            .I(N__40940));
    LocalMux I__8883 (
            .O(N__40948),
            .I(N__40940));
    InMux I__8882 (
            .O(N__40947),
            .I(N__40937));
    Span4Mux_v I__8881 (
            .O(N__40940),
            .I(N__40934));
    LocalMux I__8880 (
            .O(N__40937),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__8879 (
            .O(N__40934),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__8878 (
            .O(N__40929),
            .I(N__40926));
    LocalMux I__8877 (
            .O(N__40926),
            .I(N__40922));
    InMux I__8876 (
            .O(N__40925),
            .I(N__40918));
    Span4Mux_h I__8875 (
            .O(N__40922),
            .I(N__40915));
    InMux I__8874 (
            .O(N__40921),
            .I(N__40912));
    LocalMux I__8873 (
            .O(N__40918),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__8872 (
            .O(N__40915),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    LocalMux I__8871 (
            .O(N__40912),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    CascadeMux I__8870 (
            .O(N__40905),
            .I(N__40902));
    InMux I__8869 (
            .O(N__40902),
            .I(N__40899));
    LocalMux I__8868 (
            .O(N__40899),
            .I(N__40896));
    Odrv4 I__8867 (
            .O(N__40896),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    InMux I__8866 (
            .O(N__40893),
            .I(N__40890));
    LocalMux I__8865 (
            .O(N__40890),
            .I(N__40887));
    Span4Mux_h I__8864 (
            .O(N__40887),
            .I(N__40884));
    Odrv4 I__8863 (
            .O(N__40884),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__8862 (
            .O(N__40881),
            .I(N__40878));
    LocalMux I__8861 (
            .O(N__40878),
            .I(N__40875));
    Span4Mux_h I__8860 (
            .O(N__40875),
            .I(N__40872));
    Odrv4 I__8859 (
            .O(N__40872),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    InMux I__8858 (
            .O(N__40869),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__8857 (
            .O(N__40866),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__8856 (
            .O(N__40863),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__8855 (
            .O(N__40860),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__8854 (
            .O(N__40857),
            .I(bfn_17_10_0_));
    InMux I__8853 (
            .O(N__40854),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__8852 (
            .O(N__40851),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__8851 (
            .O(N__40848),
            .I(N__40841));
    InMux I__8850 (
            .O(N__40847),
            .I(N__40841));
    InMux I__8849 (
            .O(N__40846),
            .I(N__40838));
    LocalMux I__8848 (
            .O(N__40841),
            .I(N__40835));
    LocalMux I__8847 (
            .O(N__40838),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv12 I__8846 (
            .O(N__40835),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__8845 (
            .O(N__40830),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    CascadeMux I__8844 (
            .O(N__40827),
            .I(N__40824));
    InMux I__8843 (
            .O(N__40824),
            .I(N__40817));
    InMux I__8842 (
            .O(N__40823),
            .I(N__40817));
    InMux I__8841 (
            .O(N__40822),
            .I(N__40814));
    LocalMux I__8840 (
            .O(N__40817),
            .I(N__40811));
    LocalMux I__8839 (
            .O(N__40814),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv12 I__8838 (
            .O(N__40811),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__8837 (
            .O(N__40806),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__8836 (
            .O(N__40803),
            .I(N__40799));
    InMux I__8835 (
            .O(N__40802),
            .I(N__40796));
    LocalMux I__8834 (
            .O(N__40799),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__8833 (
            .O(N__40796),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__8832 (
            .O(N__40791),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__8831 (
            .O(N__40788),
            .I(N__40784));
    InMux I__8830 (
            .O(N__40787),
            .I(N__40781));
    LocalMux I__8829 (
            .O(N__40784),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__8828 (
            .O(N__40781),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__8827 (
            .O(N__40776),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__8826 (
            .O(N__40773),
            .I(N__40769));
    InMux I__8825 (
            .O(N__40772),
            .I(N__40766));
    LocalMux I__8824 (
            .O(N__40769),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__8823 (
            .O(N__40766),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__8822 (
            .O(N__40761),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__8821 (
            .O(N__40758),
            .I(N__40754));
    InMux I__8820 (
            .O(N__40757),
            .I(N__40751));
    LocalMux I__8819 (
            .O(N__40754),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__8818 (
            .O(N__40751),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__8817 (
            .O(N__40746),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__8816 (
            .O(N__40743),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__8815 (
            .O(N__40740),
            .I(bfn_17_9_0_));
    CascadeMux I__8814 (
            .O(N__40737),
            .I(N__40734));
    InMux I__8813 (
            .O(N__40734),
            .I(N__40728));
    InMux I__8812 (
            .O(N__40733),
            .I(N__40728));
    LocalMux I__8811 (
            .O(N__40728),
            .I(N__40724));
    InMux I__8810 (
            .O(N__40727),
            .I(N__40721));
    Span4Mux_v I__8809 (
            .O(N__40724),
            .I(N__40718));
    LocalMux I__8808 (
            .O(N__40721),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__8807 (
            .O(N__40718),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__8806 (
            .O(N__40713),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__8805 (
            .O(N__40710),
            .I(N__40704));
    InMux I__8804 (
            .O(N__40709),
            .I(N__40704));
    LocalMux I__8803 (
            .O(N__40704),
            .I(N__40700));
    InMux I__8802 (
            .O(N__40703),
            .I(N__40697));
    Span4Mux_h I__8801 (
            .O(N__40700),
            .I(N__40694));
    LocalMux I__8800 (
            .O(N__40697),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__8799 (
            .O(N__40694),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__8798 (
            .O(N__40689),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__8797 (
            .O(N__40686),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__8796 (
            .O(N__40683),
            .I(N__40679));
    InMux I__8795 (
            .O(N__40682),
            .I(N__40676));
    LocalMux I__8794 (
            .O(N__40679),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__8793 (
            .O(N__40676),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__8792 (
            .O(N__40671),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__8791 (
            .O(N__40668),
            .I(N__40664));
    InMux I__8790 (
            .O(N__40667),
            .I(N__40661));
    LocalMux I__8789 (
            .O(N__40664),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__8788 (
            .O(N__40661),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__8787 (
            .O(N__40656),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__8786 (
            .O(N__40653),
            .I(N__40649));
    InMux I__8785 (
            .O(N__40652),
            .I(N__40646));
    LocalMux I__8784 (
            .O(N__40649),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__8783 (
            .O(N__40646),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__8782 (
            .O(N__40641),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__8781 (
            .O(N__40638),
            .I(N__40634));
    InMux I__8780 (
            .O(N__40637),
            .I(N__40631));
    LocalMux I__8779 (
            .O(N__40634),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__8778 (
            .O(N__40631),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__8777 (
            .O(N__40626),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__8776 (
            .O(N__40623),
            .I(N__40619));
    InMux I__8775 (
            .O(N__40622),
            .I(N__40616));
    LocalMux I__8774 (
            .O(N__40619),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__8773 (
            .O(N__40616),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__8772 (
            .O(N__40611),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__8771 (
            .O(N__40608),
            .I(N__40604));
    InMux I__8770 (
            .O(N__40607),
            .I(N__40601));
    LocalMux I__8769 (
            .O(N__40604),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__8768 (
            .O(N__40601),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__8767 (
            .O(N__40596),
            .I(bfn_17_8_0_));
    InMux I__8766 (
            .O(N__40593),
            .I(N__40589));
    InMux I__8765 (
            .O(N__40592),
            .I(N__40586));
    LocalMux I__8764 (
            .O(N__40589),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__8763 (
            .O(N__40586),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__8762 (
            .O(N__40581),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__8761 (
            .O(N__40578),
            .I(N__40574));
    InMux I__8760 (
            .O(N__40577),
            .I(N__40571));
    LocalMux I__8759 (
            .O(N__40574),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__8758 (
            .O(N__40571),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__8757 (
            .O(N__40566),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    CascadeMux I__8756 (
            .O(N__40563),
            .I(N__40559));
    CascadeMux I__8755 (
            .O(N__40562),
            .I(N__40556));
    InMux I__8754 (
            .O(N__40559),
            .I(N__40553));
    InMux I__8753 (
            .O(N__40556),
            .I(N__40549));
    LocalMux I__8752 (
            .O(N__40553),
            .I(N__40545));
    InMux I__8751 (
            .O(N__40552),
            .I(N__40542));
    LocalMux I__8750 (
            .O(N__40549),
            .I(N__40539));
    InMux I__8749 (
            .O(N__40548),
            .I(N__40536));
    Span4Mux_v I__8748 (
            .O(N__40545),
            .I(N__40533));
    LocalMux I__8747 (
            .O(N__40542),
            .I(N__40530));
    Span4Mux_h I__8746 (
            .O(N__40539),
            .I(N__40525));
    LocalMux I__8745 (
            .O(N__40536),
            .I(N__40525));
    Odrv4 I__8744 (
            .O(N__40533),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__8743 (
            .O(N__40530),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__8742 (
            .O(N__40525),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    CascadeMux I__8741 (
            .O(N__40518),
            .I(N__40515));
    InMux I__8740 (
            .O(N__40515),
            .I(N__40512));
    LocalMux I__8739 (
            .O(N__40512),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__8738 (
            .O(N__40509),
            .I(N__40506));
    InMux I__8737 (
            .O(N__40506),
            .I(N__40503));
    LocalMux I__8736 (
            .O(N__40503),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__8735 (
            .O(N__40500),
            .I(N__40497));
    LocalMux I__8734 (
            .O(N__40497),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__8733 (
            .O(N__40494),
            .I(N__40491));
    InMux I__8732 (
            .O(N__40491),
            .I(N__40488));
    LocalMux I__8731 (
            .O(N__40488),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__8730 (
            .O(N__40485),
            .I(N__40482));
    LocalMux I__8729 (
            .O(N__40482),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    InMux I__8728 (
            .O(N__40479),
            .I(N__40474));
    InMux I__8727 (
            .O(N__40478),
            .I(N__40469));
    InMux I__8726 (
            .O(N__40477),
            .I(N__40469));
    LocalMux I__8725 (
            .O(N__40474),
            .I(N__40465));
    LocalMux I__8724 (
            .O(N__40469),
            .I(N__40462));
    InMux I__8723 (
            .O(N__40468),
            .I(N__40459));
    Span4Mux_h I__8722 (
            .O(N__40465),
            .I(N__40454));
    Span4Mux_h I__8721 (
            .O(N__40462),
            .I(N__40454));
    LocalMux I__8720 (
            .O(N__40459),
            .I(N__40451));
    Span4Mux_v I__8719 (
            .O(N__40454),
            .I(N__40448));
    Span4Mux_h I__8718 (
            .O(N__40451),
            .I(N__40445));
    Odrv4 I__8717 (
            .O(N__40448),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__8716 (
            .O(N__40445),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__8715 (
            .O(N__40440),
            .I(N__40437));
    LocalMux I__8714 (
            .O(N__40437),
            .I(N__40433));
    InMux I__8713 (
            .O(N__40436),
            .I(N__40430));
    Odrv12 I__8712 (
            .O(N__40433),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    LocalMux I__8711 (
            .O(N__40430),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__8710 (
            .O(N__40425),
            .I(N__40422));
    LocalMux I__8709 (
            .O(N__40422),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    CascadeMux I__8708 (
            .O(N__40419),
            .I(N__40415));
    InMux I__8707 (
            .O(N__40418),
            .I(N__40411));
    InMux I__8706 (
            .O(N__40415),
            .I(N__40408));
    InMux I__8705 (
            .O(N__40414),
            .I(N__40405));
    LocalMux I__8704 (
            .O(N__40411),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__8703 (
            .O(N__40408),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__8702 (
            .O(N__40405),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__8701 (
            .O(N__40398),
            .I(N__40394));
    InMux I__8700 (
            .O(N__40397),
            .I(N__40391));
    LocalMux I__8699 (
            .O(N__40394),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__8698 (
            .O(N__40391),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__8697 (
            .O(N__40386),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__8696 (
            .O(N__40383),
            .I(N__40380));
    InMux I__8695 (
            .O(N__40380),
            .I(N__40377));
    LocalMux I__8694 (
            .O(N__40377),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ));
    InMux I__8693 (
            .O(N__40374),
            .I(N__40370));
    InMux I__8692 (
            .O(N__40373),
            .I(N__40367));
    LocalMux I__8691 (
            .O(N__40370),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__8690 (
            .O(N__40367),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__8689 (
            .O(N__40362),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__8688 (
            .O(N__40359),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__8687 (
            .O(N__40356),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__8686 (
            .O(N__40353),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__8685 (
            .O(N__40350),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__8684 (
            .O(N__40347),
            .I(N__40344));
    InMux I__8683 (
            .O(N__40344),
            .I(N__40341));
    LocalMux I__8682 (
            .O(N__40341),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__8681 (
            .O(N__40338),
            .I(N__40335));
    LocalMux I__8680 (
            .O(N__40335),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__8679 (
            .O(N__40332),
            .I(N__40329));
    LocalMux I__8678 (
            .O(N__40329),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__8677 (
            .O(N__40326),
            .I(N__40321));
    InMux I__8676 (
            .O(N__40325),
            .I(N__40318));
    InMux I__8675 (
            .O(N__40324),
            .I(N__40314));
    LocalMux I__8674 (
            .O(N__40321),
            .I(N__40309));
    LocalMux I__8673 (
            .O(N__40318),
            .I(N__40309));
    InMux I__8672 (
            .O(N__40317),
            .I(N__40306));
    LocalMux I__8671 (
            .O(N__40314),
            .I(N__40303));
    Span4Mux_h I__8670 (
            .O(N__40309),
            .I(N__40298));
    LocalMux I__8669 (
            .O(N__40306),
            .I(N__40298));
    Odrv12 I__8668 (
            .O(N__40303),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__8667 (
            .O(N__40298),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    CascadeMux I__8666 (
            .O(N__40293),
            .I(N__40290));
    InMux I__8665 (
            .O(N__40290),
            .I(N__40287));
    LocalMux I__8664 (
            .O(N__40287),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__8663 (
            .O(N__40284),
            .I(N__40281));
    InMux I__8662 (
            .O(N__40281),
            .I(N__40278));
    LocalMux I__8661 (
            .O(N__40278),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__8660 (
            .O(N__40275),
            .I(bfn_16_21_0_));
    InMux I__8659 (
            .O(N__40272),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__8658 (
            .O(N__40269),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__8657 (
            .O(N__40266),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__8656 (
            .O(N__40263),
            .I(N__40260));
    InMux I__8655 (
            .O(N__40260),
            .I(N__40257));
    LocalMux I__8654 (
            .O(N__40257),
            .I(N__40253));
    InMux I__8653 (
            .O(N__40256),
            .I(N__40250));
    Sp12to4 I__8652 (
            .O(N__40253),
            .I(N__40245));
    LocalMux I__8651 (
            .O(N__40250),
            .I(N__40242));
    InMux I__8650 (
            .O(N__40249),
            .I(N__40237));
    InMux I__8649 (
            .O(N__40248),
            .I(N__40237));
    Span12Mux_v I__8648 (
            .O(N__40245),
            .I(N__40234));
    Span4Mux_v I__8647 (
            .O(N__40242),
            .I(N__40229));
    LocalMux I__8646 (
            .O(N__40237),
            .I(N__40229));
    Odrv12 I__8645 (
            .O(N__40234),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__8644 (
            .O(N__40229),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__8643 (
            .O(N__40224),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__8642 (
            .O(N__40221),
            .I(N__40217));
    InMux I__8641 (
            .O(N__40220),
            .I(N__40214));
    LocalMux I__8640 (
            .O(N__40217),
            .I(N__40210));
    LocalMux I__8639 (
            .O(N__40214),
            .I(N__40207));
    InMux I__8638 (
            .O(N__40213),
            .I(N__40204));
    Span4Mux_v I__8637 (
            .O(N__40210),
            .I(N__40200));
    Span4Mux_h I__8636 (
            .O(N__40207),
            .I(N__40197));
    LocalMux I__8635 (
            .O(N__40204),
            .I(N__40194));
    InMux I__8634 (
            .O(N__40203),
            .I(N__40191));
    Odrv4 I__8633 (
            .O(N__40200),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__8632 (
            .O(N__40197),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__8631 (
            .O(N__40194),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__8630 (
            .O(N__40191),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__8629 (
            .O(N__40182),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__8628 (
            .O(N__40179),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__8627 (
            .O(N__40176),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__8626 (
            .O(N__40173),
            .I(bfn_16_22_0_));
    CascadeMux I__8625 (
            .O(N__40170),
            .I(N__40167));
    InMux I__8624 (
            .O(N__40167),
            .I(N__40163));
    CascadeMux I__8623 (
            .O(N__40166),
            .I(N__40160));
    LocalMux I__8622 (
            .O(N__40163),
            .I(N__40155));
    InMux I__8621 (
            .O(N__40160),
            .I(N__40152));
    InMux I__8620 (
            .O(N__40159),
            .I(N__40147));
    InMux I__8619 (
            .O(N__40158),
            .I(N__40147));
    Sp12to4 I__8618 (
            .O(N__40155),
            .I(N__40142));
    LocalMux I__8617 (
            .O(N__40152),
            .I(N__40142));
    LocalMux I__8616 (
            .O(N__40147),
            .I(N__40139));
    Odrv12 I__8615 (
            .O(N__40142),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__8614 (
            .O(N__40139),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__8613 (
            .O(N__40134),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__8612 (
            .O(N__40131),
            .I(bfn_16_20_0_));
    InMux I__8611 (
            .O(N__40128),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__8610 (
            .O(N__40125),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__8609 (
            .O(N__40122),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__8608 (
            .O(N__40119),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__8607 (
            .O(N__40116),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__8606 (
            .O(N__40113),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__8605 (
            .O(N__40110),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__8604 (
            .O(N__40107),
            .I(N__40104));
    LocalMux I__8603 (
            .O(N__40104),
            .I(N__40101));
    Span4Mux_v I__8602 (
            .O(N__40101),
            .I(N__40098));
    Odrv4 I__8601 (
            .O(N__40098),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__8600 (
            .O(N__40095),
            .I(N__40091));
    CascadeMux I__8599 (
            .O(N__40094),
            .I(N__40088));
    InMux I__8598 (
            .O(N__40091),
            .I(N__40085));
    InMux I__8597 (
            .O(N__40088),
            .I(N__40082));
    LocalMux I__8596 (
            .O(N__40085),
            .I(N__40075));
    LocalMux I__8595 (
            .O(N__40082),
            .I(N__40075));
    InMux I__8594 (
            .O(N__40081),
            .I(N__40072));
    InMux I__8593 (
            .O(N__40080),
            .I(N__40069));
    Span4Mux_v I__8592 (
            .O(N__40075),
            .I(N__40066));
    LocalMux I__8591 (
            .O(N__40072),
            .I(N__40063));
    LocalMux I__8590 (
            .O(N__40069),
            .I(N__40060));
    Odrv4 I__8589 (
            .O(N__40066),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv12 I__8588 (
            .O(N__40063),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__8587 (
            .O(N__40060),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__8586 (
            .O(N__40053),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__8585 (
            .O(N__40050),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__8584 (
            .O(N__40047),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__8583 (
            .O(N__40044),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__8582 (
            .O(N__40041),
            .I(N__40038));
    InMux I__8581 (
            .O(N__40038),
            .I(N__40034));
    CascadeMux I__8580 (
            .O(N__40037),
            .I(N__40031));
    LocalMux I__8579 (
            .O(N__40034),
            .I(N__40028));
    InMux I__8578 (
            .O(N__40031),
            .I(N__40024));
    Span4Mux_h I__8577 (
            .O(N__40028),
            .I(N__40021));
    InMux I__8576 (
            .O(N__40027),
            .I(N__40018));
    LocalMux I__8575 (
            .O(N__40024),
            .I(N__40015));
    Span4Mux_v I__8574 (
            .O(N__40021),
            .I(N__40012));
    LocalMux I__8573 (
            .O(N__40018),
            .I(N__40009));
    Span4Mux_v I__8572 (
            .O(N__40015),
            .I(N__40005));
    Span4Mux_h I__8571 (
            .O(N__40012),
            .I(N__40002));
    Span4Mux_v I__8570 (
            .O(N__40009),
            .I(N__39999));
    InMux I__8569 (
            .O(N__40008),
            .I(N__39996));
    Odrv4 I__8568 (
            .O(N__40005),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__8567 (
            .O(N__40002),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__8566 (
            .O(N__39999),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__8565 (
            .O(N__39996),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__8564 (
            .O(N__39987),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__8563 (
            .O(N__39984),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__8562 (
            .O(N__39981),
            .I(N__39978));
    InMux I__8561 (
            .O(N__39978),
            .I(N__39975));
    LocalMux I__8560 (
            .O(N__39975),
            .I(N__39972));
    Span4Mux_v I__8559 (
            .O(N__39972),
            .I(N__39969));
    Odrv4 I__8558 (
            .O(N__39969),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    CascadeMux I__8557 (
            .O(N__39966),
            .I(N__39963));
    InMux I__8556 (
            .O(N__39963),
            .I(N__39960));
    LocalMux I__8555 (
            .O(N__39960),
            .I(N__39957));
    Odrv12 I__8554 (
            .O(N__39957),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    CascadeMux I__8553 (
            .O(N__39954),
            .I(N__39951));
    InMux I__8552 (
            .O(N__39951),
            .I(N__39948));
    LocalMux I__8551 (
            .O(N__39948),
            .I(N__39945));
    Span4Mux_v I__8550 (
            .O(N__39945),
            .I(N__39942));
    Odrv4 I__8549 (
            .O(N__39942),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    CascadeMux I__8548 (
            .O(N__39939),
            .I(N__39936));
    InMux I__8547 (
            .O(N__39936),
            .I(N__39933));
    LocalMux I__8546 (
            .O(N__39933),
            .I(N__39930));
    Span4Mux_h I__8545 (
            .O(N__39930),
            .I(N__39927));
    Odrv4 I__8544 (
            .O(N__39927),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    CascadeMux I__8543 (
            .O(N__39924),
            .I(N__39921));
    InMux I__8542 (
            .O(N__39921),
            .I(N__39918));
    LocalMux I__8541 (
            .O(N__39918),
            .I(N__39915));
    Span4Mux_v I__8540 (
            .O(N__39915),
            .I(N__39912));
    Odrv4 I__8539 (
            .O(N__39912),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__8538 (
            .O(N__39909),
            .I(N__39906));
    LocalMux I__8537 (
            .O(N__39906),
            .I(N__39903));
    Span4Mux_v I__8536 (
            .O(N__39903),
            .I(N__39900));
    Odrv4 I__8535 (
            .O(N__39900),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    InMux I__8534 (
            .O(N__39897),
            .I(N__39894));
    LocalMux I__8533 (
            .O(N__39894),
            .I(N__39891));
    Odrv4 I__8532 (
            .O(N__39891),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ));
    CascadeMux I__8531 (
            .O(N__39888),
            .I(N__39885));
    InMux I__8530 (
            .O(N__39885),
            .I(N__39882));
    LocalMux I__8529 (
            .O(N__39882),
            .I(N__39879));
    Span4Mux_v I__8528 (
            .O(N__39879),
            .I(N__39876));
    Span4Mux_v I__8527 (
            .O(N__39876),
            .I(N__39873));
    Odrv4 I__8526 (
            .O(N__39873),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__8525 (
            .O(N__39870),
            .I(N__39867));
    LocalMux I__8524 (
            .O(N__39867),
            .I(N__39864));
    Span4Mux_v I__8523 (
            .O(N__39864),
            .I(N__39861));
    Odrv4 I__8522 (
            .O(N__39861),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__8521 (
            .O(N__39858),
            .I(N__39855));
    LocalMux I__8520 (
            .O(N__39855),
            .I(N__39852));
    Span4Mux_v I__8519 (
            .O(N__39852),
            .I(N__39849));
    Span4Mux_v I__8518 (
            .O(N__39849),
            .I(N__39846));
    Odrv4 I__8517 (
            .O(N__39846),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    CascadeMux I__8516 (
            .O(N__39843),
            .I(N__39840));
    InMux I__8515 (
            .O(N__39840),
            .I(N__39837));
    LocalMux I__8514 (
            .O(N__39837),
            .I(N__39834));
    Span4Mux_v I__8513 (
            .O(N__39834),
            .I(N__39831));
    Odrv4 I__8512 (
            .O(N__39831),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__8511 (
            .O(N__39828),
            .I(N__39825));
    LocalMux I__8510 (
            .O(N__39825),
            .I(N__39822));
    Span4Mux_v I__8509 (
            .O(N__39822),
            .I(N__39819));
    Odrv4 I__8508 (
            .O(N__39819),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__8507 (
            .O(N__39816),
            .I(N__39813));
    InMux I__8506 (
            .O(N__39813),
            .I(N__39810));
    LocalMux I__8505 (
            .O(N__39810),
            .I(N__39807));
    Span4Mux_v I__8504 (
            .O(N__39807),
            .I(N__39804));
    Odrv4 I__8503 (
            .O(N__39804),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__8502 (
            .O(N__39801),
            .I(N__39798));
    LocalMux I__8501 (
            .O(N__39798),
            .I(N__39795));
    Span4Mux_v I__8500 (
            .O(N__39795),
            .I(N__39792));
    Odrv4 I__8499 (
            .O(N__39792),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    InMux I__8498 (
            .O(N__39789),
            .I(N__39786));
    LocalMux I__8497 (
            .O(N__39786),
            .I(N__39783));
    Span4Mux_h I__8496 (
            .O(N__39783),
            .I(N__39780));
    Odrv4 I__8495 (
            .O(N__39780),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    CascadeMux I__8494 (
            .O(N__39777),
            .I(N__39774));
    InMux I__8493 (
            .O(N__39774),
            .I(N__39771));
    LocalMux I__8492 (
            .O(N__39771),
            .I(N__39768));
    Span4Mux_v I__8491 (
            .O(N__39768),
            .I(N__39765));
    Odrv4 I__8490 (
            .O(N__39765),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ));
    InMux I__8489 (
            .O(N__39762),
            .I(N__39759));
    LocalMux I__8488 (
            .O(N__39759),
            .I(N__39756));
    Span4Mux_v I__8487 (
            .O(N__39756),
            .I(N__39753));
    Odrv4 I__8486 (
            .O(N__39753),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    InMux I__8485 (
            .O(N__39750),
            .I(N__39747));
    LocalMux I__8484 (
            .O(N__39747),
            .I(N__39744));
    Span4Mux_h I__8483 (
            .O(N__39744),
            .I(N__39741));
    Odrv4 I__8482 (
            .O(N__39741),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ));
    InMux I__8481 (
            .O(N__39738),
            .I(N__39735));
    LocalMux I__8480 (
            .O(N__39735),
            .I(N__39732));
    Span4Mux_v I__8479 (
            .O(N__39732),
            .I(N__39729));
    Odrv4 I__8478 (
            .O(N__39729),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__8477 (
            .O(N__39726),
            .I(N__39723));
    LocalMux I__8476 (
            .O(N__39723),
            .I(N__39720));
    Span4Mux_v I__8475 (
            .O(N__39720),
            .I(N__39717));
    Span4Mux_v I__8474 (
            .O(N__39717),
            .I(N__39714));
    Odrv4 I__8473 (
            .O(N__39714),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__8472 (
            .O(N__39711),
            .I(N__39708));
    InMux I__8471 (
            .O(N__39708),
            .I(N__39705));
    LocalMux I__8470 (
            .O(N__39705),
            .I(N__39702));
    Span4Mux_v I__8469 (
            .O(N__39702),
            .I(N__39699));
    Odrv4 I__8468 (
            .O(N__39699),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__8467 (
            .O(N__39696),
            .I(N__39690));
    InMux I__8466 (
            .O(N__39695),
            .I(N__39685));
    InMux I__8465 (
            .O(N__39694),
            .I(N__39685));
    InMux I__8464 (
            .O(N__39693),
            .I(N__39682));
    LocalMux I__8463 (
            .O(N__39690),
            .I(N__39679));
    LocalMux I__8462 (
            .O(N__39685),
            .I(N__39676));
    LocalMux I__8461 (
            .O(N__39682),
            .I(N__39673));
    Span4Mux_h I__8460 (
            .O(N__39679),
            .I(N__39670));
    Span4Mux_v I__8459 (
            .O(N__39676),
            .I(N__39667));
    Span4Mux_v I__8458 (
            .O(N__39673),
            .I(N__39664));
    Odrv4 I__8457 (
            .O(N__39670),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__8456 (
            .O(N__39667),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__8455 (
            .O(N__39664),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__8454 (
            .O(N__39657),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8453 (
            .O(N__39654),
            .I(N__39650));
    InMux I__8452 (
            .O(N__39653),
            .I(N__39645));
    LocalMux I__8451 (
            .O(N__39650),
            .I(N__39642));
    InMux I__8450 (
            .O(N__39649),
            .I(N__39639));
    InMux I__8449 (
            .O(N__39648),
            .I(N__39636));
    LocalMux I__8448 (
            .O(N__39645),
            .I(N__39633));
    Span4Mux_v I__8447 (
            .O(N__39642),
            .I(N__39626));
    LocalMux I__8446 (
            .O(N__39639),
            .I(N__39626));
    LocalMux I__8445 (
            .O(N__39636),
            .I(N__39626));
    Span4Mux_v I__8444 (
            .O(N__39633),
            .I(N__39623));
    Span4Mux_h I__8443 (
            .O(N__39626),
            .I(N__39620));
    Odrv4 I__8442 (
            .O(N__39623),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    Odrv4 I__8441 (
            .O(N__39620),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__8440 (
            .O(N__39615),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__8439 (
            .O(N__39612),
            .I(N__39607));
    InMux I__8438 (
            .O(N__39611),
            .I(N__39604));
    CascadeMux I__8437 (
            .O(N__39610),
            .I(N__39601));
    LocalMux I__8436 (
            .O(N__39607),
            .I(N__39595));
    LocalMux I__8435 (
            .O(N__39604),
            .I(N__39595));
    InMux I__8434 (
            .O(N__39601),
            .I(N__39592));
    InMux I__8433 (
            .O(N__39600),
            .I(N__39589));
    Span4Mux_v I__8432 (
            .O(N__39595),
            .I(N__39584));
    LocalMux I__8431 (
            .O(N__39592),
            .I(N__39584));
    LocalMux I__8430 (
            .O(N__39589),
            .I(N__39581));
    Span4Mux_h I__8429 (
            .O(N__39584),
            .I(N__39578));
    Odrv12 I__8428 (
            .O(N__39581),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__8427 (
            .O(N__39578),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__8426 (
            .O(N__39573),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8425 (
            .O(N__39570),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__8424 (
            .O(N__39567),
            .I(N__39564));
    LocalMux I__8423 (
            .O(N__39564),
            .I(N__39558));
    InMux I__8422 (
            .O(N__39563),
            .I(N__39555));
    InMux I__8421 (
            .O(N__39562),
            .I(N__39550));
    InMux I__8420 (
            .O(N__39561),
            .I(N__39550));
    Span4Mux_v I__8419 (
            .O(N__39558),
            .I(N__39543));
    LocalMux I__8418 (
            .O(N__39555),
            .I(N__39543));
    LocalMux I__8417 (
            .O(N__39550),
            .I(N__39543));
    Span4Mux_h I__8416 (
            .O(N__39543),
            .I(N__39540));
    Odrv4 I__8415 (
            .O(N__39540),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    CascadeMux I__8414 (
            .O(N__39537),
            .I(N__39534));
    InMux I__8413 (
            .O(N__39534),
            .I(N__39529));
    InMux I__8412 (
            .O(N__39533),
            .I(N__39526));
    CascadeMux I__8411 (
            .O(N__39532),
            .I(N__39522));
    LocalMux I__8410 (
            .O(N__39529),
            .I(N__39517));
    LocalMux I__8409 (
            .O(N__39526),
            .I(N__39517));
    InMux I__8408 (
            .O(N__39525),
            .I(N__39512));
    InMux I__8407 (
            .O(N__39522),
            .I(N__39512));
    Span4Mux_v I__8406 (
            .O(N__39517),
            .I(N__39507));
    LocalMux I__8405 (
            .O(N__39512),
            .I(N__39507));
    Odrv4 I__8404 (
            .O(N__39507),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__8403 (
            .O(N__39504),
            .I(N__39501));
    LocalMux I__8402 (
            .O(N__39501),
            .I(N__39498));
    Span4Mux_h I__8401 (
            .O(N__39498),
            .I(N__39495));
    Odrv4 I__8400 (
            .O(N__39495),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ));
    CascadeMux I__8399 (
            .O(N__39492),
            .I(N__39489));
    InMux I__8398 (
            .O(N__39489),
            .I(N__39486));
    LocalMux I__8397 (
            .O(N__39486),
            .I(N__39483));
    Span4Mux_v I__8396 (
            .O(N__39483),
            .I(N__39480));
    Odrv4 I__8395 (
            .O(N__39480),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    InMux I__8394 (
            .O(N__39477),
            .I(N__39474));
    LocalMux I__8393 (
            .O(N__39474),
            .I(N__39471));
    Span4Mux_v I__8392 (
            .O(N__39471),
            .I(N__39468));
    Odrv4 I__8391 (
            .O(N__39468),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    InMux I__8390 (
            .O(N__39465),
            .I(N__39461));
    InMux I__8389 (
            .O(N__39464),
            .I(N__39457));
    LocalMux I__8388 (
            .O(N__39461),
            .I(N__39454));
    InMux I__8387 (
            .O(N__39460),
            .I(N__39451));
    LocalMux I__8386 (
            .O(N__39457),
            .I(N__39447));
    Span4Mux_h I__8385 (
            .O(N__39454),
            .I(N__39442));
    LocalMux I__8384 (
            .O(N__39451),
            .I(N__39442));
    InMux I__8383 (
            .O(N__39450),
            .I(N__39439));
    Span4Mux_v I__8382 (
            .O(N__39447),
            .I(N__39436));
    Odrv4 I__8381 (
            .O(N__39442),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    LocalMux I__8380 (
            .O(N__39439),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__8379 (
            .O(N__39436),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__8378 (
            .O(N__39429),
            .I(bfn_16_12_0_));
    InMux I__8377 (
            .O(N__39426),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__8376 (
            .O(N__39423),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__8375 (
            .O(N__39420),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__8374 (
            .O(N__39417),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__8373 (
            .O(N__39414),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__8372 (
            .O(N__39411),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__8371 (
            .O(N__39408),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__8370 (
            .O(N__39405),
            .I(bfn_16_13_0_));
    InMux I__8369 (
            .O(N__39402),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__8368 (
            .O(N__39399),
            .I(bfn_16_11_0_));
    InMux I__8367 (
            .O(N__39396),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__8366 (
            .O(N__39393),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__8365 (
            .O(N__39390),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__8364 (
            .O(N__39387),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__8363 (
            .O(N__39384),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__8362 (
            .O(N__39381),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__8361 (
            .O(N__39378),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__8360 (
            .O(N__39375),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    InMux I__8359 (
            .O(N__39372),
            .I(N__39365));
    InMux I__8358 (
            .O(N__39371),
            .I(N__39365));
    InMux I__8357 (
            .O(N__39370),
            .I(N__39362));
    LocalMux I__8356 (
            .O(N__39365),
            .I(N__39357));
    LocalMux I__8355 (
            .O(N__39362),
            .I(N__39357));
    Odrv12 I__8354 (
            .O(N__39357),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__8353 (
            .O(N__39354),
            .I(N__39349));
    InMux I__8352 (
            .O(N__39353),
            .I(N__39346));
    InMux I__8351 (
            .O(N__39352),
            .I(N__39343));
    LocalMux I__8350 (
            .O(N__39349),
            .I(N__39338));
    LocalMux I__8349 (
            .O(N__39346),
            .I(N__39338));
    LocalMux I__8348 (
            .O(N__39343),
            .I(N__39334));
    Span4Mux_v I__8347 (
            .O(N__39338),
            .I(N__39331));
    InMux I__8346 (
            .O(N__39337),
            .I(N__39328));
    Odrv4 I__8345 (
            .O(N__39334),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__8344 (
            .O(N__39331),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__8343 (
            .O(N__39328),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__8342 (
            .O(N__39321),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__8341 (
            .O(N__39318),
            .I(N__39310));
    InMux I__8340 (
            .O(N__39317),
            .I(N__39310));
    InMux I__8339 (
            .O(N__39316),
            .I(N__39307));
    InMux I__8338 (
            .O(N__39315),
            .I(N__39304));
    LocalMux I__8337 (
            .O(N__39310),
            .I(N__39301));
    LocalMux I__8336 (
            .O(N__39307),
            .I(N__39298));
    LocalMux I__8335 (
            .O(N__39304),
            .I(N__39295));
    Span4Mux_h I__8334 (
            .O(N__39301),
            .I(N__39292));
    Span4Mux_v I__8333 (
            .O(N__39298),
            .I(N__39289));
    Odrv4 I__8332 (
            .O(N__39295),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__8331 (
            .O(N__39292),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__8330 (
            .O(N__39289),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__8329 (
            .O(N__39282),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__8328 (
            .O(N__39279),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__8327 (
            .O(N__39276),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__8326 (
            .O(N__39273),
            .I(N__39269));
    InMux I__8325 (
            .O(N__39272),
            .I(N__39265));
    LocalMux I__8324 (
            .O(N__39269),
            .I(N__39261));
    InMux I__8323 (
            .O(N__39268),
            .I(N__39258));
    LocalMux I__8322 (
            .O(N__39265),
            .I(N__39255));
    InMux I__8321 (
            .O(N__39264),
            .I(N__39252));
    Span4Mux_v I__8320 (
            .O(N__39261),
            .I(N__39247));
    LocalMux I__8319 (
            .O(N__39258),
            .I(N__39247));
    Span4Mux_h I__8318 (
            .O(N__39255),
            .I(N__39240));
    LocalMux I__8317 (
            .O(N__39252),
            .I(N__39240));
    Span4Mux_h I__8316 (
            .O(N__39247),
            .I(N__39240));
    Span4Mux_v I__8315 (
            .O(N__39240),
            .I(N__39237));
    Odrv4 I__8314 (
            .O(N__39237),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__8313 (
            .O(N__39234),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__8312 (
            .O(N__39231),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__8311 (
            .O(N__39228),
            .I(N__39225));
    LocalMux I__8310 (
            .O(N__39225),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__8309 (
            .O(N__39222),
            .I(N__39219));
    LocalMux I__8308 (
            .O(N__39219),
            .I(N__39216));
    Span4Mux_v I__8307 (
            .O(N__39216),
            .I(N__39213));
    Odrv4 I__8306 (
            .O(N__39213),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    CascadeMux I__8305 (
            .O(N__39210),
            .I(N__39207));
    InMux I__8304 (
            .O(N__39207),
            .I(N__39204));
    LocalMux I__8303 (
            .O(N__39204),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    InMux I__8302 (
            .O(N__39201),
            .I(N__39198));
    LocalMux I__8301 (
            .O(N__39198),
            .I(N__39195));
    Span4Mux_v I__8300 (
            .O(N__39195),
            .I(N__39192));
    Span4Mux_h I__8299 (
            .O(N__39192),
            .I(N__39189));
    Odrv4 I__8298 (
            .O(N__39189),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    CascadeMux I__8297 (
            .O(N__39186),
            .I(N__39183));
    InMux I__8296 (
            .O(N__39183),
            .I(N__39180));
    LocalMux I__8295 (
            .O(N__39180),
            .I(N__39177));
    Span4Mux_v I__8294 (
            .O(N__39177),
            .I(N__39174));
    Odrv4 I__8293 (
            .O(N__39174),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    InMux I__8292 (
            .O(N__39171),
            .I(N__39168));
    LocalMux I__8291 (
            .O(N__39168),
            .I(N__39165));
    Odrv4 I__8290 (
            .O(N__39165),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    CascadeMux I__8289 (
            .O(N__39162),
            .I(N__39159));
    InMux I__8288 (
            .O(N__39159),
            .I(N__39156));
    LocalMux I__8287 (
            .O(N__39156),
            .I(N__39153));
    Span4Mux_h I__8286 (
            .O(N__39153),
            .I(N__39150));
    Odrv4 I__8285 (
            .O(N__39150),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    CascadeMux I__8284 (
            .O(N__39147),
            .I(N__39144));
    InMux I__8283 (
            .O(N__39144),
            .I(N__39141));
    LocalMux I__8282 (
            .O(N__39141),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__8281 (
            .O(N__39138),
            .I(N__39135));
    LocalMux I__8280 (
            .O(N__39135),
            .I(N__39132));
    Span4Mux_v I__8279 (
            .O(N__39132),
            .I(N__39129));
    Span4Mux_h I__8278 (
            .O(N__39129),
            .I(N__39126));
    Odrv4 I__8277 (
            .O(N__39126),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__8276 (
            .O(N__39123),
            .I(N__39120));
    InMux I__8275 (
            .O(N__39120),
            .I(N__39117));
    LocalMux I__8274 (
            .O(N__39117),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__8273 (
            .O(N__39114),
            .I(N__39111));
    InMux I__8272 (
            .O(N__39111),
            .I(N__39108));
    LocalMux I__8271 (
            .O(N__39108),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__8270 (
            .O(N__39105),
            .I(N__39102));
    InMux I__8269 (
            .O(N__39102),
            .I(N__39099));
    LocalMux I__8268 (
            .O(N__39099),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__8267 (
            .O(N__39096),
            .I(N__39093));
    LocalMux I__8266 (
            .O(N__39093),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__8265 (
            .O(N__39090),
            .I(N__39087));
    InMux I__8264 (
            .O(N__39087),
            .I(N__39084));
    LocalMux I__8263 (
            .O(N__39084),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__8262 (
            .O(N__39081),
            .I(N__39078));
    InMux I__8261 (
            .O(N__39078),
            .I(N__39075));
    LocalMux I__8260 (
            .O(N__39075),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__8259 (
            .O(N__39072),
            .I(N__39069));
    InMux I__8258 (
            .O(N__39069),
            .I(N__39066));
    LocalMux I__8257 (
            .O(N__39066),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__8256 (
            .O(N__39063),
            .I(N__39052));
    InMux I__8255 (
            .O(N__39062),
            .I(N__39052));
    InMux I__8254 (
            .O(N__39061),
            .I(N__39052));
    InMux I__8253 (
            .O(N__39060),
            .I(N__39047));
    InMux I__8252 (
            .O(N__39059),
            .I(N__39047));
    LocalMux I__8251 (
            .O(N__39052),
            .I(N__39044));
    LocalMux I__8250 (
            .O(N__39047),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__8249 (
            .O(N__39044),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    CascadeMux I__8248 (
            .O(N__39039),
            .I(N__39036));
    InMux I__8247 (
            .O(N__39036),
            .I(N__39030));
    InMux I__8246 (
            .O(N__39035),
            .I(N__39030));
    LocalMux I__8245 (
            .O(N__39030),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__8244 (
            .O(N__39027),
            .I(N__39023));
    CascadeMux I__8243 (
            .O(N__39026),
            .I(N__39020));
    InMux I__8242 (
            .O(N__39023),
            .I(N__39013));
    InMux I__8241 (
            .O(N__39020),
            .I(N__39013));
    InMux I__8240 (
            .O(N__39019),
            .I(N__39008));
    InMux I__8239 (
            .O(N__39018),
            .I(N__39008));
    LocalMux I__8238 (
            .O(N__39013),
            .I(N__39005));
    LocalMux I__8237 (
            .O(N__39008),
            .I(N__39002));
    Span4Mux_h I__8236 (
            .O(N__39005),
            .I(N__38998));
    Span4Mux_h I__8235 (
            .O(N__39002),
            .I(N__38995));
    InMux I__8234 (
            .O(N__39001),
            .I(N__38992));
    Odrv4 I__8233 (
            .O(N__38998),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__8232 (
            .O(N__38995),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__8231 (
            .O(N__38992),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    InMux I__8230 (
            .O(N__38985),
            .I(N__38981));
    InMux I__8229 (
            .O(N__38984),
            .I(N__38976));
    LocalMux I__8228 (
            .O(N__38981),
            .I(N__38973));
    InMux I__8227 (
            .O(N__38980),
            .I(N__38970));
    CascadeMux I__8226 (
            .O(N__38979),
            .I(N__38967));
    LocalMux I__8225 (
            .O(N__38976),
            .I(N__38960));
    Span4Mux_v I__8224 (
            .O(N__38973),
            .I(N__38960));
    LocalMux I__8223 (
            .O(N__38970),
            .I(N__38960));
    InMux I__8222 (
            .O(N__38967),
            .I(N__38957));
    Span4Mux_h I__8221 (
            .O(N__38960),
            .I(N__38954));
    LocalMux I__8220 (
            .O(N__38957),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__8219 (
            .O(N__38954),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    CascadeMux I__8218 (
            .O(N__38949),
            .I(N__38946));
    InMux I__8217 (
            .O(N__38946),
            .I(N__38943));
    LocalMux I__8216 (
            .O(N__38943),
            .I(N__38940));
    Odrv4 I__8215 (
            .O(N__38940),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__8214 (
            .O(N__38937),
            .I(N__38934));
    LocalMux I__8213 (
            .O(N__38934),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__8212 (
            .O(N__38931),
            .I(N__38928));
    InMux I__8211 (
            .O(N__38928),
            .I(N__38925));
    LocalMux I__8210 (
            .O(N__38925),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__8209 (
            .O(N__38922),
            .I(N__38919));
    LocalMux I__8208 (
            .O(N__38919),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__8207 (
            .O(N__38916),
            .I(N__38913));
    InMux I__8206 (
            .O(N__38913),
            .I(N__38910));
    LocalMux I__8205 (
            .O(N__38910),
            .I(N__38907));
    Odrv4 I__8204 (
            .O(N__38907),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__8203 (
            .O(N__38904),
            .I(N__38901));
    LocalMux I__8202 (
            .O(N__38901),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__8201 (
            .O(N__38898),
            .I(N__38895));
    InMux I__8200 (
            .O(N__38895),
            .I(N__38892));
    LocalMux I__8199 (
            .O(N__38892),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__8198 (
            .O(N__38889),
            .I(N__38886));
    LocalMux I__8197 (
            .O(N__38886),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__8196 (
            .O(N__38883),
            .I(N__38880));
    InMux I__8195 (
            .O(N__38880),
            .I(N__38877));
    LocalMux I__8194 (
            .O(N__38877),
            .I(N__38874));
    Odrv4 I__8193 (
            .O(N__38874),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__8192 (
            .O(N__38871),
            .I(N__38868));
    InMux I__8191 (
            .O(N__38868),
            .I(N__38865));
    LocalMux I__8190 (
            .O(N__38865),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__8189 (
            .O(N__38862),
            .I(N__38845));
    InMux I__8188 (
            .O(N__38861),
            .I(N__38838));
    InMux I__8187 (
            .O(N__38860),
            .I(N__38838));
    InMux I__8186 (
            .O(N__38859),
            .I(N__38838));
    InMux I__8185 (
            .O(N__38858),
            .I(N__38829));
    InMux I__8184 (
            .O(N__38857),
            .I(N__38829));
    InMux I__8183 (
            .O(N__38856),
            .I(N__38829));
    InMux I__8182 (
            .O(N__38855),
            .I(N__38829));
    CascadeMux I__8181 (
            .O(N__38854),
            .I(N__38825));
    CascadeMux I__8180 (
            .O(N__38853),
            .I(N__38821));
    CascadeMux I__8179 (
            .O(N__38852),
            .I(N__38817));
    CascadeMux I__8178 (
            .O(N__38851),
            .I(N__38812));
    CascadeMux I__8177 (
            .O(N__38850),
            .I(N__38808));
    CascadeMux I__8176 (
            .O(N__38849),
            .I(N__38804));
    InMux I__8175 (
            .O(N__38848),
            .I(N__38800));
    LocalMux I__8174 (
            .O(N__38845),
            .I(N__38793));
    LocalMux I__8173 (
            .O(N__38838),
            .I(N__38793));
    LocalMux I__8172 (
            .O(N__38829),
            .I(N__38793));
    InMux I__8171 (
            .O(N__38828),
            .I(N__38778));
    InMux I__8170 (
            .O(N__38825),
            .I(N__38778));
    InMux I__8169 (
            .O(N__38824),
            .I(N__38778));
    InMux I__8168 (
            .O(N__38821),
            .I(N__38778));
    InMux I__8167 (
            .O(N__38820),
            .I(N__38778));
    InMux I__8166 (
            .O(N__38817),
            .I(N__38778));
    InMux I__8165 (
            .O(N__38816),
            .I(N__38778));
    InMux I__8164 (
            .O(N__38815),
            .I(N__38763));
    InMux I__8163 (
            .O(N__38812),
            .I(N__38763));
    InMux I__8162 (
            .O(N__38811),
            .I(N__38763));
    InMux I__8161 (
            .O(N__38808),
            .I(N__38763));
    InMux I__8160 (
            .O(N__38807),
            .I(N__38763));
    InMux I__8159 (
            .O(N__38804),
            .I(N__38763));
    InMux I__8158 (
            .O(N__38803),
            .I(N__38763));
    LocalMux I__8157 (
            .O(N__38800),
            .I(N__38750));
    Span4Mux_v I__8156 (
            .O(N__38793),
            .I(N__38743));
    LocalMux I__8155 (
            .O(N__38778),
            .I(N__38740));
    LocalMux I__8154 (
            .O(N__38763),
            .I(N__38737));
    CascadeMux I__8153 (
            .O(N__38762),
            .I(N__38733));
    CascadeMux I__8152 (
            .O(N__38761),
            .I(N__38729));
    CascadeMux I__8151 (
            .O(N__38760),
            .I(N__38725));
    CascadeMux I__8150 (
            .O(N__38759),
            .I(N__38721));
    InMux I__8149 (
            .O(N__38758),
            .I(N__38718));
    InMux I__8148 (
            .O(N__38757),
            .I(N__38713));
    InMux I__8147 (
            .O(N__38756),
            .I(N__38713));
    InMux I__8146 (
            .O(N__38755),
            .I(N__38710));
    InMux I__8145 (
            .O(N__38754),
            .I(N__38703));
    InMux I__8144 (
            .O(N__38753),
            .I(N__38700));
    Span4Mux_s1_h I__8143 (
            .O(N__38750),
            .I(N__38697));
    CascadeMux I__8142 (
            .O(N__38749),
            .I(N__38694));
    CascadeMux I__8141 (
            .O(N__38748),
            .I(N__38690));
    CascadeMux I__8140 (
            .O(N__38747),
            .I(N__38686));
    CascadeMux I__8139 (
            .O(N__38746),
            .I(N__38682));
    Sp12to4 I__8138 (
            .O(N__38743),
            .I(N__38667));
    Span4Mux_v I__8137 (
            .O(N__38740),
            .I(N__38662));
    Span4Mux_v I__8136 (
            .O(N__38737),
            .I(N__38662));
    InMux I__8135 (
            .O(N__38736),
            .I(N__38645));
    InMux I__8134 (
            .O(N__38733),
            .I(N__38645));
    InMux I__8133 (
            .O(N__38732),
            .I(N__38645));
    InMux I__8132 (
            .O(N__38729),
            .I(N__38645));
    InMux I__8131 (
            .O(N__38728),
            .I(N__38645));
    InMux I__8130 (
            .O(N__38725),
            .I(N__38645));
    InMux I__8129 (
            .O(N__38724),
            .I(N__38645));
    InMux I__8128 (
            .O(N__38721),
            .I(N__38645));
    LocalMux I__8127 (
            .O(N__38718),
            .I(N__38638));
    LocalMux I__8126 (
            .O(N__38713),
            .I(N__38638));
    LocalMux I__8125 (
            .O(N__38710),
            .I(N__38638));
    InMux I__8124 (
            .O(N__38709),
            .I(N__38635));
    InMux I__8123 (
            .O(N__38708),
            .I(N__38630));
    InMux I__8122 (
            .O(N__38707),
            .I(N__38630));
    InMux I__8121 (
            .O(N__38706),
            .I(N__38627));
    LocalMux I__8120 (
            .O(N__38703),
            .I(N__38622));
    LocalMux I__8119 (
            .O(N__38700),
            .I(N__38622));
    Sp12to4 I__8118 (
            .O(N__38697),
            .I(N__38619));
    InMux I__8117 (
            .O(N__38694),
            .I(N__38602));
    InMux I__8116 (
            .O(N__38693),
            .I(N__38602));
    InMux I__8115 (
            .O(N__38690),
            .I(N__38602));
    InMux I__8114 (
            .O(N__38689),
            .I(N__38602));
    InMux I__8113 (
            .O(N__38686),
            .I(N__38602));
    InMux I__8112 (
            .O(N__38685),
            .I(N__38602));
    InMux I__8111 (
            .O(N__38682),
            .I(N__38602));
    InMux I__8110 (
            .O(N__38681),
            .I(N__38602));
    InMux I__8109 (
            .O(N__38680),
            .I(N__38599));
    InMux I__8108 (
            .O(N__38679),
            .I(N__38596));
    InMux I__8107 (
            .O(N__38678),
            .I(N__38593));
    InMux I__8106 (
            .O(N__38677),
            .I(N__38590));
    InMux I__8105 (
            .O(N__38676),
            .I(N__38583));
    InMux I__8104 (
            .O(N__38675),
            .I(N__38583));
    InMux I__8103 (
            .O(N__38674),
            .I(N__38583));
    InMux I__8102 (
            .O(N__38673),
            .I(N__38574));
    InMux I__8101 (
            .O(N__38672),
            .I(N__38574));
    InMux I__8100 (
            .O(N__38671),
            .I(N__38574));
    InMux I__8099 (
            .O(N__38670),
            .I(N__38574));
    Span12Mux_s8_h I__8098 (
            .O(N__38667),
            .I(N__38565));
    Sp12to4 I__8097 (
            .O(N__38662),
            .I(N__38565));
    LocalMux I__8096 (
            .O(N__38645),
            .I(N__38565));
    Span12Mux_s9_v I__8095 (
            .O(N__38638),
            .I(N__38556));
    LocalMux I__8094 (
            .O(N__38635),
            .I(N__38556));
    LocalMux I__8093 (
            .O(N__38630),
            .I(N__38556));
    LocalMux I__8092 (
            .O(N__38627),
            .I(N__38556));
    Span4Mux_v I__8091 (
            .O(N__38622),
            .I(N__38553));
    Span12Mux_s8_v I__8090 (
            .O(N__38619),
            .I(N__38548));
    LocalMux I__8089 (
            .O(N__38602),
            .I(N__38548));
    LocalMux I__8088 (
            .O(N__38599),
            .I(N__38535));
    LocalMux I__8087 (
            .O(N__38596),
            .I(N__38535));
    LocalMux I__8086 (
            .O(N__38593),
            .I(N__38535));
    LocalMux I__8085 (
            .O(N__38590),
            .I(N__38535));
    LocalMux I__8084 (
            .O(N__38583),
            .I(N__38535));
    LocalMux I__8083 (
            .O(N__38574),
            .I(N__38535));
    CascadeMux I__8082 (
            .O(N__38573),
            .I(N__38532));
    CascadeMux I__8081 (
            .O(N__38572),
            .I(N__38528));
    Span12Mux_h I__8080 (
            .O(N__38565),
            .I(N__38525));
    Span12Mux_v I__8079 (
            .O(N__38556),
            .I(N__38516));
    Sp12to4 I__8078 (
            .O(N__38553),
            .I(N__38516));
    Span12Mux_h I__8077 (
            .O(N__38548),
            .I(N__38516));
    Span12Mux_s8_v I__8076 (
            .O(N__38535),
            .I(N__38516));
    InMux I__8075 (
            .O(N__38532),
            .I(N__38509));
    InMux I__8074 (
            .O(N__38531),
            .I(N__38509));
    InMux I__8073 (
            .O(N__38528),
            .I(N__38509));
    Odrv12 I__8072 (
            .O(N__38525),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__8071 (
            .O(N__38516),
            .I(CONSTANT_ONE_NET));
    LocalMux I__8070 (
            .O(N__38509),
            .I(CONSTANT_ONE_NET));
    InMux I__8069 (
            .O(N__38502),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    CascadeMux I__8068 (
            .O(N__38499),
            .I(N__38486));
    InMux I__8067 (
            .O(N__38498),
            .I(N__38480));
    InMux I__8066 (
            .O(N__38497),
            .I(N__38480));
    InMux I__8065 (
            .O(N__38496),
            .I(N__38476));
    InMux I__8064 (
            .O(N__38495),
            .I(N__38471));
    InMux I__8063 (
            .O(N__38494),
            .I(N__38471));
    InMux I__8062 (
            .O(N__38493),
            .I(N__38468));
    CascadeMux I__8061 (
            .O(N__38492),
            .I(N__38464));
    InMux I__8060 (
            .O(N__38491),
            .I(N__38449));
    InMux I__8059 (
            .O(N__38490),
            .I(N__38449));
    InMux I__8058 (
            .O(N__38489),
            .I(N__38446));
    InMux I__8057 (
            .O(N__38486),
            .I(N__38443));
    InMux I__8056 (
            .O(N__38485),
            .I(N__38439));
    LocalMux I__8055 (
            .O(N__38480),
            .I(N__38436));
    InMux I__8054 (
            .O(N__38479),
            .I(N__38433));
    LocalMux I__8053 (
            .O(N__38476),
            .I(N__38419));
    LocalMux I__8052 (
            .O(N__38471),
            .I(N__38419));
    LocalMux I__8051 (
            .O(N__38468),
            .I(N__38419));
    InMux I__8050 (
            .O(N__38467),
            .I(N__38406));
    InMux I__8049 (
            .O(N__38464),
            .I(N__38406));
    InMux I__8048 (
            .O(N__38463),
            .I(N__38406));
    InMux I__8047 (
            .O(N__38462),
            .I(N__38406));
    InMux I__8046 (
            .O(N__38461),
            .I(N__38406));
    InMux I__8045 (
            .O(N__38460),
            .I(N__38406));
    InMux I__8044 (
            .O(N__38459),
            .I(N__38393));
    InMux I__8043 (
            .O(N__38458),
            .I(N__38393));
    InMux I__8042 (
            .O(N__38457),
            .I(N__38393));
    InMux I__8041 (
            .O(N__38456),
            .I(N__38393));
    InMux I__8040 (
            .O(N__38455),
            .I(N__38393));
    InMux I__8039 (
            .O(N__38454),
            .I(N__38393));
    LocalMux I__8038 (
            .O(N__38449),
            .I(N__38388));
    LocalMux I__8037 (
            .O(N__38446),
            .I(N__38388));
    LocalMux I__8036 (
            .O(N__38443),
            .I(N__38385));
    InMux I__8035 (
            .O(N__38442),
            .I(N__38382));
    LocalMux I__8034 (
            .O(N__38439),
            .I(N__38379));
    Span4Mux_v I__8033 (
            .O(N__38436),
            .I(N__38374));
    LocalMux I__8032 (
            .O(N__38433),
            .I(N__38374));
    InMux I__8031 (
            .O(N__38432),
            .I(N__38365));
    InMux I__8030 (
            .O(N__38431),
            .I(N__38365));
    InMux I__8029 (
            .O(N__38430),
            .I(N__38365));
    InMux I__8028 (
            .O(N__38429),
            .I(N__38365));
    InMux I__8027 (
            .O(N__38428),
            .I(N__38358));
    InMux I__8026 (
            .O(N__38427),
            .I(N__38358));
    InMux I__8025 (
            .O(N__38426),
            .I(N__38358));
    Sp12to4 I__8024 (
            .O(N__38419),
            .I(N__38349));
    LocalMux I__8023 (
            .O(N__38406),
            .I(N__38349));
    LocalMux I__8022 (
            .O(N__38393),
            .I(N__38349));
    Sp12to4 I__8021 (
            .O(N__38388),
            .I(N__38349));
    Span4Mux_v I__8020 (
            .O(N__38385),
            .I(N__38340));
    LocalMux I__8019 (
            .O(N__38382),
            .I(N__38340));
    Span4Mux_h I__8018 (
            .O(N__38379),
            .I(N__38340));
    Span4Mux_h I__8017 (
            .O(N__38374),
            .I(N__38340));
    LocalMux I__8016 (
            .O(N__38365),
            .I(N__38335));
    LocalMux I__8015 (
            .O(N__38358),
            .I(N__38335));
    Span12Mux_v I__8014 (
            .O(N__38349),
            .I(N__38332));
    Sp12to4 I__8013 (
            .O(N__38340),
            .I(N__38327));
    Span12Mux_v I__8012 (
            .O(N__38335),
            .I(N__38327));
    Odrv12 I__8011 (
            .O(N__38332),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv12 I__8010 (
            .O(N__38327),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    CascadeMux I__8009 (
            .O(N__38322),
            .I(N__38317));
    InMux I__8008 (
            .O(N__38321),
            .I(N__38313));
    InMux I__8007 (
            .O(N__38320),
            .I(N__38310));
    InMux I__8006 (
            .O(N__38317),
            .I(N__38307));
    InMux I__8005 (
            .O(N__38316),
            .I(N__38304));
    LocalMux I__8004 (
            .O(N__38313),
            .I(N__38297));
    LocalMux I__8003 (
            .O(N__38310),
            .I(N__38297));
    LocalMux I__8002 (
            .O(N__38307),
            .I(N__38297));
    LocalMux I__8001 (
            .O(N__38304),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__8000 (
            .O(N__38297),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__7999 (
            .O(N__38292),
            .I(N__38288));
    InMux I__7998 (
            .O(N__38291),
            .I(N__38285));
    LocalMux I__7997 (
            .O(N__38288),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    LocalMux I__7996 (
            .O(N__38285),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    CascadeMux I__7995 (
            .O(N__38280),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__7994 (
            .O(N__38277),
            .I(N__38273));
    InMux I__7993 (
            .O(N__38276),
            .I(N__38268));
    InMux I__7992 (
            .O(N__38273),
            .I(N__38265));
    InMux I__7991 (
            .O(N__38272),
            .I(N__38260));
    InMux I__7990 (
            .O(N__38271),
            .I(N__38260));
    LocalMux I__7989 (
            .O(N__38268),
            .I(N__38257));
    LocalMux I__7988 (
            .O(N__38265),
            .I(N__38254));
    LocalMux I__7987 (
            .O(N__38260),
            .I(N__38250));
    Span4Mux_v I__7986 (
            .O(N__38257),
            .I(N__38244));
    Span4Mux_h I__7985 (
            .O(N__38254),
            .I(N__38244));
    InMux I__7984 (
            .O(N__38253),
            .I(N__38241));
    Span12Mux_v I__7983 (
            .O(N__38250),
            .I(N__38238));
    InMux I__7982 (
            .O(N__38249),
            .I(N__38235));
    Odrv4 I__7981 (
            .O(N__38244),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__7980 (
            .O(N__38241),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv12 I__7979 (
            .O(N__38238),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__7978 (
            .O(N__38235),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__7977 (
            .O(N__38226),
            .I(N__38223));
    LocalMux I__7976 (
            .O(N__38223),
            .I(N__38220));
    Odrv4 I__7975 (
            .O(N__38220),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    CascadeMux I__7974 (
            .O(N__38217),
            .I(N__38214));
    InMux I__7973 (
            .O(N__38214),
            .I(N__38211));
    LocalMux I__7972 (
            .O(N__38211),
            .I(N__38208));
    Odrv4 I__7971 (
            .O(N__38208),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    InMux I__7970 (
            .O(N__38205),
            .I(N__38202));
    LocalMux I__7969 (
            .O(N__38202),
            .I(N__38199));
    Odrv4 I__7968 (
            .O(N__38199),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    CascadeMux I__7967 (
            .O(N__38196),
            .I(N__38193));
    InMux I__7966 (
            .O(N__38193),
            .I(N__38190));
    LocalMux I__7965 (
            .O(N__38190),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    CascadeMux I__7964 (
            .O(N__38187),
            .I(N__38184));
    InMux I__7963 (
            .O(N__38184),
            .I(N__38181));
    LocalMux I__7962 (
            .O(N__38181),
            .I(N__38178));
    Odrv4 I__7961 (
            .O(N__38178),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    CascadeMux I__7960 (
            .O(N__38175),
            .I(N__38172));
    InMux I__7959 (
            .O(N__38172),
            .I(N__38169));
    LocalMux I__7958 (
            .O(N__38169),
            .I(N__38166));
    Odrv4 I__7957 (
            .O(N__38166),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__7956 (
            .O(N__38163),
            .I(N__38160));
    LocalMux I__7955 (
            .O(N__38160),
            .I(N__38157));
    Odrv12 I__7954 (
            .O(N__38157),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__7953 (
            .O(N__38154),
            .I(N__38151));
    LocalMux I__7952 (
            .O(N__38151),
            .I(N__38148));
    Odrv4 I__7951 (
            .O(N__38148),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__7950 (
            .O(N__38145),
            .I(N__38142));
    LocalMux I__7949 (
            .O(N__38142),
            .I(N__38139));
    Span4Mux_h I__7948 (
            .O(N__38139),
            .I(N__38136));
    Odrv4 I__7947 (
            .O(N__38136),
            .I(\current_shift_inst.control_input_axb_4 ));
    CascadeMux I__7946 (
            .O(N__38133),
            .I(N__38130));
    InMux I__7945 (
            .O(N__38130),
            .I(N__38127));
    LocalMux I__7944 (
            .O(N__38127),
            .I(N__38124));
    Odrv4 I__7943 (
            .O(N__38124),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__7942 (
            .O(N__38121),
            .I(N__38118));
    LocalMux I__7941 (
            .O(N__38118),
            .I(N__38115));
    Odrv4 I__7940 (
            .O(N__38115),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__7939 (
            .O(N__38112),
            .I(N__38109));
    LocalMux I__7938 (
            .O(N__38109),
            .I(N__38106));
    Span4Mux_h I__7937 (
            .O(N__38106),
            .I(N__38103));
    Odrv4 I__7936 (
            .O(N__38103),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__7935 (
            .O(N__38100),
            .I(N__38097));
    LocalMux I__7934 (
            .O(N__38097),
            .I(N__38094));
    Span4Mux_h I__7933 (
            .O(N__38094),
            .I(N__38091));
    Odrv4 I__7932 (
            .O(N__38091),
            .I(\current_shift_inst.control_input_axb_7 ));
    CascadeMux I__7931 (
            .O(N__38088),
            .I(N__38085));
    InMux I__7930 (
            .O(N__38085),
            .I(N__38082));
    LocalMux I__7929 (
            .O(N__38082),
            .I(N__38079));
    Odrv4 I__7928 (
            .O(N__38079),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__7927 (
            .O(N__38076),
            .I(N__38073));
    LocalMux I__7926 (
            .O(N__38073),
            .I(N__38070));
    Odrv4 I__7925 (
            .O(N__38070),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    CascadeMux I__7924 (
            .O(N__38067),
            .I(N__38064));
    InMux I__7923 (
            .O(N__38064),
            .I(N__38061));
    LocalMux I__7922 (
            .O(N__38061),
            .I(N__38058));
    Span4Mux_h I__7921 (
            .O(N__38058),
            .I(N__38055));
    Odrv4 I__7920 (
            .O(N__38055),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__7919 (
            .O(N__38052),
            .I(N__38049));
    LocalMux I__7918 (
            .O(N__38049),
            .I(N__38046));
    Span4Mux_v I__7917 (
            .O(N__38046),
            .I(N__38043));
    Odrv4 I__7916 (
            .O(N__38043),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__7915 (
            .O(N__38040),
            .I(N__38037));
    LocalMux I__7914 (
            .O(N__38037),
            .I(N__38034));
    Odrv4 I__7913 (
            .O(N__38034),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__7912 (
            .O(N__38031),
            .I(N__38028));
    LocalMux I__7911 (
            .O(N__38028),
            .I(N__38025));
    Odrv4 I__7910 (
            .O(N__38025),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__7909 (
            .O(N__38022),
            .I(N__38019));
    LocalMux I__7908 (
            .O(N__38019),
            .I(N__38016));
    Span4Mux_h I__7907 (
            .O(N__38016),
            .I(N__38013));
    Odrv4 I__7906 (
            .O(N__38013),
            .I(\current_shift_inst.control_input_axb_3 ));
    CascadeMux I__7905 (
            .O(N__38010),
            .I(N__38007));
    InMux I__7904 (
            .O(N__38007),
            .I(N__38004));
    LocalMux I__7903 (
            .O(N__38004),
            .I(N__38001));
    Odrv4 I__7902 (
            .O(N__38001),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    InMux I__7901 (
            .O(N__37998),
            .I(N__37995));
    LocalMux I__7900 (
            .O(N__37995),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__7899 (
            .O(N__37992),
            .I(N__37989));
    LocalMux I__7898 (
            .O(N__37989),
            .I(N__37986));
    Odrv4 I__7897 (
            .O(N__37986),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    CascadeMux I__7896 (
            .O(N__37983),
            .I(N__37980));
    InMux I__7895 (
            .O(N__37980),
            .I(N__37977));
    LocalMux I__7894 (
            .O(N__37977),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    CascadeMux I__7893 (
            .O(N__37974),
            .I(N__37971));
    InMux I__7892 (
            .O(N__37971),
            .I(N__37968));
    LocalMux I__7891 (
            .O(N__37968),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__7890 (
            .O(N__37965),
            .I(N__37962));
    LocalMux I__7889 (
            .O(N__37962),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    CascadeMux I__7888 (
            .O(N__37959),
            .I(N__37956));
    InMux I__7887 (
            .O(N__37956),
            .I(N__37953));
    LocalMux I__7886 (
            .O(N__37953),
            .I(N__37950));
    Span4Mux_h I__7885 (
            .O(N__37950),
            .I(N__37947));
    Odrv4 I__7884 (
            .O(N__37947),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    CascadeMux I__7883 (
            .O(N__37944),
            .I(N__37941));
    InMux I__7882 (
            .O(N__37941),
            .I(N__37938));
    LocalMux I__7881 (
            .O(N__37938),
            .I(N__37935));
    Odrv4 I__7880 (
            .O(N__37935),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    CascadeMux I__7879 (
            .O(N__37932),
            .I(N__37929));
    InMux I__7878 (
            .O(N__37929),
            .I(N__37926));
    LocalMux I__7877 (
            .O(N__37926),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    InMux I__7876 (
            .O(N__37923),
            .I(N__37920));
    LocalMux I__7875 (
            .O(N__37920),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    InMux I__7874 (
            .O(N__37917),
            .I(N__37914));
    LocalMux I__7873 (
            .O(N__37914),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__7872 (
            .O(N__37911),
            .I(N__37908));
    LocalMux I__7871 (
            .O(N__37908),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__7870 (
            .O(N__37905),
            .I(N__37902));
    LocalMux I__7869 (
            .O(N__37902),
            .I(N__37897));
    InMux I__7868 (
            .O(N__37901),
            .I(N__37894));
    InMux I__7867 (
            .O(N__37900),
            .I(N__37891));
    Span4Mux_v I__7866 (
            .O(N__37897),
            .I(N__37886));
    LocalMux I__7865 (
            .O(N__37894),
            .I(N__37886));
    LocalMux I__7864 (
            .O(N__37891),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    Odrv4 I__7863 (
            .O(N__37886),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    InMux I__7862 (
            .O(N__37881),
            .I(N__37878));
    LocalMux I__7861 (
            .O(N__37878),
            .I(N__37875));
    Span4Mux_h I__7860 (
            .O(N__37875),
            .I(N__37872));
    Span4Mux_v I__7859 (
            .O(N__37872),
            .I(N__37869));
    Odrv4 I__7858 (
            .O(N__37869),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__7857 (
            .O(N__37866),
            .I(N__37863));
    LocalMux I__7856 (
            .O(N__37863),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__7855 (
            .O(N__37860),
            .I(N__37857));
    LocalMux I__7854 (
            .O(N__37857),
            .I(N__37854));
    Span4Mux_h I__7853 (
            .O(N__37854),
            .I(N__37851));
    Odrv4 I__7852 (
            .O(N__37851),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__7851 (
            .O(N__37848),
            .I(N__37845));
    LocalMux I__7850 (
            .O(N__37845),
            .I(\current_shift_inst.un38_control_input_0_s0_3 ));
    InMux I__7849 (
            .O(N__37842),
            .I(N__37839));
    LocalMux I__7848 (
            .O(N__37839),
            .I(N__37836));
    Span4Mux_h I__7847 (
            .O(N__37836),
            .I(N__37833));
    Odrv4 I__7846 (
            .O(N__37833),
            .I(\current_shift_inst.un38_control_input_0_s1_3 ));
    InMux I__7845 (
            .O(N__37830),
            .I(N__37826));
    InMux I__7844 (
            .O(N__37829),
            .I(N__37823));
    LocalMux I__7843 (
            .O(N__37826),
            .I(N__37818));
    LocalMux I__7842 (
            .O(N__37823),
            .I(N__37818));
    Odrv12 I__7841 (
            .O(N__37818),
            .I(\current_shift_inst.control_input_axb_0 ));
    InMux I__7840 (
            .O(N__37815),
            .I(N__37812));
    LocalMux I__7839 (
            .O(N__37812),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ));
    CascadeMux I__7838 (
            .O(N__37809),
            .I(N__37806));
    InMux I__7837 (
            .O(N__37806),
            .I(N__37803));
    LocalMux I__7836 (
            .O(N__37803),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    InMux I__7835 (
            .O(N__37800),
            .I(N__37797));
    LocalMux I__7834 (
            .O(N__37797),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    CascadeMux I__7833 (
            .O(N__37794),
            .I(N__37791));
    InMux I__7832 (
            .O(N__37791),
            .I(N__37788));
    LocalMux I__7831 (
            .O(N__37788),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    InMux I__7830 (
            .O(N__37785),
            .I(N__37782));
    LocalMux I__7829 (
            .O(N__37782),
            .I(N__37779));
    Odrv12 I__7828 (
            .O(N__37779),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    CascadeMux I__7827 (
            .O(N__37776),
            .I(N__37773));
    InMux I__7826 (
            .O(N__37773),
            .I(N__37770));
    LocalMux I__7825 (
            .O(N__37770),
            .I(N__37767));
    Span4Mux_v I__7824 (
            .O(N__37767),
            .I(N__37764));
    Span4Mux_h I__7823 (
            .O(N__37764),
            .I(N__37761));
    Odrv4 I__7822 (
            .O(N__37761),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    CascadeMux I__7821 (
            .O(N__37758),
            .I(N__37754));
    InMux I__7820 (
            .O(N__37757),
            .I(N__37748));
    InMux I__7819 (
            .O(N__37754),
            .I(N__37748));
    InMux I__7818 (
            .O(N__37753),
            .I(N__37745));
    LocalMux I__7817 (
            .O(N__37748),
            .I(N__37742));
    LocalMux I__7816 (
            .O(N__37745),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__7815 (
            .O(N__37742),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    CascadeMux I__7814 (
            .O(N__37737),
            .I(N__37733));
    InMux I__7813 (
            .O(N__37736),
            .I(N__37727));
    InMux I__7812 (
            .O(N__37733),
            .I(N__37727));
    InMux I__7811 (
            .O(N__37732),
            .I(N__37724));
    LocalMux I__7810 (
            .O(N__37727),
            .I(N__37721));
    LocalMux I__7809 (
            .O(N__37724),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__7808 (
            .O(N__37721),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__7807 (
            .O(N__37716),
            .I(N__37713));
    LocalMux I__7806 (
            .O(N__37713),
            .I(N__37710));
    Span4Mux_h I__7805 (
            .O(N__37710),
            .I(N__37707));
    Odrv4 I__7804 (
            .O(N__37707),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    InMux I__7803 (
            .O(N__37704),
            .I(N__37698));
    InMux I__7802 (
            .O(N__37703),
            .I(N__37698));
    LocalMux I__7801 (
            .O(N__37698),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    CascadeMux I__7800 (
            .O(N__37695),
            .I(elapsed_time_ns_1_RNI03DN9_0_22_cascade_));
    InMux I__7799 (
            .O(N__37692),
            .I(N__37686));
    InMux I__7798 (
            .O(N__37691),
            .I(N__37686));
    LocalMux I__7797 (
            .O(N__37686),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    InMux I__7796 (
            .O(N__37683),
            .I(N__37680));
    LocalMux I__7795 (
            .O(N__37680),
            .I(N__37676));
    InMux I__7794 (
            .O(N__37679),
            .I(N__37672));
    Span4Mux_h I__7793 (
            .O(N__37676),
            .I(N__37669));
    InMux I__7792 (
            .O(N__37675),
            .I(N__37666));
    LocalMux I__7791 (
            .O(N__37672),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    Odrv4 I__7790 (
            .O(N__37669),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    LocalMux I__7789 (
            .O(N__37666),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    InMux I__7788 (
            .O(N__37659),
            .I(N__37656));
    LocalMux I__7787 (
            .O(N__37656),
            .I(N__37653));
    Span4Mux_h I__7786 (
            .O(N__37653),
            .I(N__37650));
    Span4Mux_v I__7785 (
            .O(N__37650),
            .I(N__37647));
    Odrv4 I__7784 (
            .O(N__37647),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    CEMux I__7783 (
            .O(N__37644),
            .I(N__37635));
    CEMux I__7782 (
            .O(N__37643),
            .I(N__37631));
    CEMux I__7781 (
            .O(N__37642),
            .I(N__37616));
    CEMux I__7780 (
            .O(N__37641),
            .I(N__37613));
    CEMux I__7779 (
            .O(N__37640),
            .I(N__37604));
    CEMux I__7778 (
            .O(N__37639),
            .I(N__37601));
    CEMux I__7777 (
            .O(N__37638),
            .I(N__37598));
    LocalMux I__7776 (
            .O(N__37635),
            .I(N__37594));
    CEMux I__7775 (
            .O(N__37634),
            .I(N__37591));
    LocalMux I__7774 (
            .O(N__37631),
            .I(N__37580));
    CEMux I__7773 (
            .O(N__37630),
            .I(N__37577));
    InMux I__7772 (
            .O(N__37629),
            .I(N__37568));
    InMux I__7771 (
            .O(N__37628),
            .I(N__37568));
    InMux I__7770 (
            .O(N__37627),
            .I(N__37568));
    InMux I__7769 (
            .O(N__37626),
            .I(N__37568));
    InMux I__7768 (
            .O(N__37625),
            .I(N__37559));
    InMux I__7767 (
            .O(N__37624),
            .I(N__37559));
    InMux I__7766 (
            .O(N__37623),
            .I(N__37559));
    InMux I__7765 (
            .O(N__37622),
            .I(N__37559));
    InMux I__7764 (
            .O(N__37621),
            .I(N__37548));
    InMux I__7763 (
            .O(N__37620),
            .I(N__37548));
    InMux I__7762 (
            .O(N__37619),
            .I(N__37548));
    LocalMux I__7761 (
            .O(N__37616),
            .I(N__37543));
    LocalMux I__7760 (
            .O(N__37613),
            .I(N__37543));
    InMux I__7759 (
            .O(N__37612),
            .I(N__37534));
    InMux I__7758 (
            .O(N__37611),
            .I(N__37534));
    InMux I__7757 (
            .O(N__37610),
            .I(N__37534));
    InMux I__7756 (
            .O(N__37609),
            .I(N__37534));
    CEMux I__7755 (
            .O(N__37608),
            .I(N__37531));
    CEMux I__7754 (
            .O(N__37607),
            .I(N__37528));
    LocalMux I__7753 (
            .O(N__37604),
            .I(N__37525));
    LocalMux I__7752 (
            .O(N__37601),
            .I(N__37520));
    LocalMux I__7751 (
            .O(N__37598),
            .I(N__37520));
    CEMux I__7750 (
            .O(N__37597),
            .I(N__37515));
    Span4Mux_v I__7749 (
            .O(N__37594),
            .I(N__37510));
    LocalMux I__7748 (
            .O(N__37591),
            .I(N__37510));
    InMux I__7747 (
            .O(N__37590),
            .I(N__37503));
    InMux I__7746 (
            .O(N__37589),
            .I(N__37496));
    InMux I__7745 (
            .O(N__37588),
            .I(N__37496));
    InMux I__7744 (
            .O(N__37587),
            .I(N__37496));
    InMux I__7743 (
            .O(N__37586),
            .I(N__37487));
    InMux I__7742 (
            .O(N__37585),
            .I(N__37487));
    InMux I__7741 (
            .O(N__37584),
            .I(N__37487));
    InMux I__7740 (
            .O(N__37583),
            .I(N__37487));
    Span4Mux_v I__7739 (
            .O(N__37580),
            .I(N__37478));
    LocalMux I__7738 (
            .O(N__37577),
            .I(N__37478));
    LocalMux I__7737 (
            .O(N__37568),
            .I(N__37478));
    LocalMux I__7736 (
            .O(N__37559),
            .I(N__37478));
    InMux I__7735 (
            .O(N__37558),
            .I(N__37469));
    InMux I__7734 (
            .O(N__37557),
            .I(N__37469));
    InMux I__7733 (
            .O(N__37556),
            .I(N__37469));
    InMux I__7732 (
            .O(N__37555),
            .I(N__37469));
    LocalMux I__7731 (
            .O(N__37548),
            .I(N__37460));
    Span4Mux_v I__7730 (
            .O(N__37543),
            .I(N__37460));
    LocalMux I__7729 (
            .O(N__37534),
            .I(N__37460));
    LocalMux I__7728 (
            .O(N__37531),
            .I(N__37460));
    LocalMux I__7727 (
            .O(N__37528),
            .I(N__37457));
    Span4Mux_h I__7726 (
            .O(N__37525),
            .I(N__37454));
    Span4Mux_v I__7725 (
            .O(N__37520),
            .I(N__37451));
    CEMux I__7724 (
            .O(N__37519),
            .I(N__37448));
    CEMux I__7723 (
            .O(N__37518),
            .I(N__37445));
    LocalMux I__7722 (
            .O(N__37515),
            .I(N__37442));
    Span4Mux_v I__7721 (
            .O(N__37510),
            .I(N__37439));
    InMux I__7720 (
            .O(N__37509),
            .I(N__37430));
    InMux I__7719 (
            .O(N__37508),
            .I(N__37430));
    InMux I__7718 (
            .O(N__37507),
            .I(N__37430));
    InMux I__7717 (
            .O(N__37506),
            .I(N__37430));
    LocalMux I__7716 (
            .O(N__37503),
            .I(N__37427));
    LocalMux I__7715 (
            .O(N__37496),
            .I(N__37416));
    LocalMux I__7714 (
            .O(N__37487),
            .I(N__37416));
    Span4Mux_v I__7713 (
            .O(N__37478),
            .I(N__37416));
    LocalMux I__7712 (
            .O(N__37469),
            .I(N__37416));
    Span4Mux_v I__7711 (
            .O(N__37460),
            .I(N__37416));
    Span4Mux_v I__7710 (
            .O(N__37457),
            .I(N__37409));
    Span4Mux_v I__7709 (
            .O(N__37454),
            .I(N__37409));
    Span4Mux_v I__7708 (
            .O(N__37451),
            .I(N__37409));
    LocalMux I__7707 (
            .O(N__37448),
            .I(N__37404));
    LocalMux I__7706 (
            .O(N__37445),
            .I(N__37404));
    Span4Mux_h I__7705 (
            .O(N__37442),
            .I(N__37397));
    Span4Mux_h I__7704 (
            .O(N__37439),
            .I(N__37397));
    LocalMux I__7703 (
            .O(N__37430),
            .I(N__37397));
    Span4Mux_v I__7702 (
            .O(N__37427),
            .I(N__37392));
    Span4Mux_v I__7701 (
            .O(N__37416),
            .I(N__37392));
    Span4Mux_v I__7700 (
            .O(N__37409),
            .I(N__37389));
    Odrv12 I__7699 (
            .O(N__37404),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__7698 (
            .O(N__37397),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__7697 (
            .O(N__37392),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__7696 (
            .O(N__37389),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    CascadeMux I__7695 (
            .O(N__37380),
            .I(N__37377));
    InMux I__7694 (
            .O(N__37377),
            .I(N__37374));
    LocalMux I__7693 (
            .O(N__37374),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__7692 (
            .O(N__37371),
            .I(N__37368));
    LocalMux I__7691 (
            .O(N__37368),
            .I(\current_shift_inst.un38_control_input_0_s0_4 ));
    InMux I__7690 (
            .O(N__37365),
            .I(N__37362));
    LocalMux I__7689 (
            .O(N__37362),
            .I(N__37359));
    Span4Mux_v I__7688 (
            .O(N__37359),
            .I(N__37356));
    Odrv4 I__7687 (
            .O(N__37356),
            .I(\current_shift_inst.un38_control_input_0_s1_4 ));
    InMux I__7686 (
            .O(N__37353),
            .I(N__37350));
    LocalMux I__7685 (
            .O(N__37350),
            .I(N__37347));
    Span4Mux_h I__7684 (
            .O(N__37347),
            .I(N__37344));
    Odrv4 I__7683 (
            .O(N__37344),
            .I(\current_shift_inst.control_input_axb_1 ));
    CascadeMux I__7682 (
            .O(N__37341),
            .I(elapsed_time_ns_1_RNI57CN9_0_18_cascade_));
    InMux I__7681 (
            .O(N__37338),
            .I(N__37332));
    InMux I__7680 (
            .O(N__37337),
            .I(N__37332));
    LocalMux I__7679 (
            .O(N__37332),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__7678 (
            .O(N__37329),
            .I(N__37324));
    InMux I__7677 (
            .O(N__37328),
            .I(N__37319));
    InMux I__7676 (
            .O(N__37327),
            .I(N__37319));
    LocalMux I__7675 (
            .O(N__37324),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__7674 (
            .O(N__37319),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__7673 (
            .O(N__37314),
            .I(N__37310));
    CascadeMux I__7672 (
            .O(N__37313),
            .I(N__37307));
    InMux I__7671 (
            .O(N__37310),
            .I(N__37302));
    InMux I__7670 (
            .O(N__37307),
            .I(N__37302));
    LocalMux I__7669 (
            .O(N__37302),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__7668 (
            .O(N__37299),
            .I(N__37294));
    InMux I__7667 (
            .O(N__37298),
            .I(N__37289));
    InMux I__7666 (
            .O(N__37297),
            .I(N__37289));
    LocalMux I__7665 (
            .O(N__37294),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__7664 (
            .O(N__37289),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__7663 (
            .O(N__37284),
            .I(N__37281));
    LocalMux I__7662 (
            .O(N__37281),
            .I(N__37278));
    Odrv4 I__7661 (
            .O(N__37278),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    InMux I__7660 (
            .O(N__37275),
            .I(N__37272));
    LocalMux I__7659 (
            .O(N__37272),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ));
    InMux I__7658 (
            .O(N__37269),
            .I(N__37266));
    LocalMux I__7657 (
            .O(N__37266),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    InMux I__7656 (
            .O(N__37263),
            .I(N__37259));
    InMux I__7655 (
            .O(N__37262),
            .I(N__37255));
    LocalMux I__7654 (
            .O(N__37259),
            .I(N__37252));
    InMux I__7653 (
            .O(N__37258),
            .I(N__37249));
    LocalMux I__7652 (
            .O(N__37255),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    Odrv4 I__7651 (
            .O(N__37252),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    LocalMux I__7650 (
            .O(N__37249),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    InMux I__7649 (
            .O(N__37242),
            .I(N__37238));
    InMux I__7648 (
            .O(N__37241),
            .I(N__37235));
    LocalMux I__7647 (
            .O(N__37238),
            .I(N__37232));
    LocalMux I__7646 (
            .O(N__37235),
            .I(N__37229));
    Span4Mux_h I__7645 (
            .O(N__37232),
            .I(N__37226));
    Odrv4 I__7644 (
            .O(N__37229),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    Odrv4 I__7643 (
            .O(N__37226),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    InMux I__7642 (
            .O(N__37221),
            .I(N__37217));
    InMux I__7641 (
            .O(N__37220),
            .I(N__37214));
    LocalMux I__7640 (
            .O(N__37217),
            .I(N__37211));
    LocalMux I__7639 (
            .O(N__37214),
            .I(N__37208));
    Span4Mux_v I__7638 (
            .O(N__37211),
            .I(N__37205));
    Odrv4 I__7637 (
            .O(N__37208),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    Odrv4 I__7636 (
            .O(N__37205),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    InMux I__7635 (
            .O(N__37200),
            .I(N__37195));
    InMux I__7634 (
            .O(N__37199),
            .I(N__37192));
    InMux I__7633 (
            .O(N__37198),
            .I(N__37189));
    LocalMux I__7632 (
            .O(N__37195),
            .I(N__37184));
    LocalMux I__7631 (
            .O(N__37192),
            .I(N__37184));
    LocalMux I__7630 (
            .O(N__37189),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__7629 (
            .O(N__37184),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__7628 (
            .O(N__37179),
            .I(N__37174));
    InMux I__7627 (
            .O(N__37178),
            .I(N__37169));
    InMux I__7626 (
            .O(N__37177),
            .I(N__37169));
    LocalMux I__7625 (
            .O(N__37174),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__7624 (
            .O(N__37169),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    CascadeMux I__7623 (
            .O(N__37164),
            .I(N__37160));
    InMux I__7622 (
            .O(N__37163),
            .I(N__37156));
    InMux I__7621 (
            .O(N__37160),
            .I(N__37151));
    InMux I__7620 (
            .O(N__37159),
            .I(N__37151));
    LocalMux I__7619 (
            .O(N__37156),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    LocalMux I__7618 (
            .O(N__37151),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__7617 (
            .O(N__37146),
            .I(N__37143));
    LocalMux I__7616 (
            .O(N__37143),
            .I(N__37140));
    Span4Mux_h I__7615 (
            .O(N__37140),
            .I(N__37137));
    Odrv4 I__7614 (
            .O(N__37137),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    CascadeMux I__7613 (
            .O(N__37134),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21_cascade_));
    CascadeMux I__7612 (
            .O(N__37131),
            .I(N__37127));
    InMux I__7611 (
            .O(N__37130),
            .I(N__37122));
    InMux I__7610 (
            .O(N__37127),
            .I(N__37122));
    LocalMux I__7609 (
            .O(N__37122),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    CascadeMux I__7608 (
            .O(N__37119),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_));
    InMux I__7607 (
            .O(N__37116),
            .I(N__37110));
    InMux I__7606 (
            .O(N__37115),
            .I(N__37110));
    LocalMux I__7605 (
            .O(N__37110),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    InMux I__7604 (
            .O(N__37107),
            .I(N__37104));
    LocalMux I__7603 (
            .O(N__37104),
            .I(N__37101));
    Span4Mux_h I__7602 (
            .O(N__37101),
            .I(N__37098));
    Odrv4 I__7601 (
            .O(N__37098),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__7600 (
            .O(N__37095),
            .I(N__37092));
    LocalMux I__7599 (
            .O(N__37092),
            .I(N__37089));
    Span4Mux_v I__7598 (
            .O(N__37089),
            .I(N__37086));
    Odrv4 I__7597 (
            .O(N__37086),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__7596 (
            .O(N__37083),
            .I(N__37080));
    InMux I__7595 (
            .O(N__37080),
            .I(N__37077));
    LocalMux I__7594 (
            .O(N__37077),
            .I(N__37074));
    Odrv12 I__7593 (
            .O(N__37074),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    CascadeMux I__7592 (
            .O(N__37071),
            .I(elapsed_time_ns_1_RNI35CN9_0_16_cascade_));
    CascadeMux I__7591 (
            .O(N__37068),
            .I(N__37064));
    InMux I__7590 (
            .O(N__37067),
            .I(N__37059));
    InMux I__7589 (
            .O(N__37064),
            .I(N__37059));
    LocalMux I__7588 (
            .O(N__37059),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__7587 (
            .O(N__37056),
            .I(N__37053));
    InMux I__7586 (
            .O(N__37053),
            .I(N__37047));
    InMux I__7585 (
            .O(N__37052),
            .I(N__37047));
    LocalMux I__7584 (
            .O(N__37047),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__7583 (
            .O(N__37044),
            .I(N__37041));
    LocalMux I__7582 (
            .O(N__37041),
            .I(N__37037));
    InMux I__7581 (
            .O(N__37040),
            .I(N__37034));
    Odrv4 I__7580 (
            .O(N__37037),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__7579 (
            .O(N__37034),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    CascadeMux I__7578 (
            .O(N__37029),
            .I(N__37026));
    InMux I__7577 (
            .O(N__37026),
            .I(N__37023));
    LocalMux I__7576 (
            .O(N__37023),
            .I(N__37020));
    Span4Mux_h I__7575 (
            .O(N__37020),
            .I(N__37017));
    Odrv4 I__7574 (
            .O(N__37017),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    CascadeMux I__7573 (
            .O(N__37014),
            .I(N__37007));
    InMux I__7572 (
            .O(N__37013),
            .I(N__37004));
    InMux I__7571 (
            .O(N__37012),
            .I(N__36997));
    InMux I__7570 (
            .O(N__37011),
            .I(N__36997));
    InMux I__7569 (
            .O(N__37010),
            .I(N__36997));
    InMux I__7568 (
            .O(N__37007),
            .I(N__36994));
    LocalMux I__7567 (
            .O(N__37004),
            .I(N__36991));
    LocalMux I__7566 (
            .O(N__36997),
            .I(N__36988));
    LocalMux I__7565 (
            .O(N__36994),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__7564 (
            .O(N__36991),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__7563 (
            .O(N__36988),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__7562 (
            .O(N__36981),
            .I(N__36975));
    InMux I__7561 (
            .O(N__36980),
            .I(N__36972));
    InMux I__7560 (
            .O(N__36979),
            .I(N__36967));
    InMux I__7559 (
            .O(N__36978),
            .I(N__36967));
    LocalMux I__7558 (
            .O(N__36975),
            .I(N__36964));
    LocalMux I__7557 (
            .O(N__36972),
            .I(N__36961));
    LocalMux I__7556 (
            .O(N__36967),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__7555 (
            .O(N__36964),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__7554 (
            .O(N__36961),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__7553 (
            .O(N__36954),
            .I(N__36950));
    InMux I__7552 (
            .O(N__36953),
            .I(N__36945));
    InMux I__7551 (
            .O(N__36950),
            .I(N__36945));
    LocalMux I__7550 (
            .O(N__36945),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    CascadeMux I__7549 (
            .O(N__36942),
            .I(elapsed_time_ns_1_RNI13CN9_0_14_cascade_));
    InMux I__7548 (
            .O(N__36939),
            .I(N__36936));
    LocalMux I__7547 (
            .O(N__36936),
            .I(N__36933));
    Span4Mux_h I__7546 (
            .O(N__36933),
            .I(N__36930));
    Odrv4 I__7545 (
            .O(N__36930),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__7544 (
            .O(N__36927),
            .I(N__36924));
    InMux I__7543 (
            .O(N__36924),
            .I(N__36921));
    LocalMux I__7542 (
            .O(N__36921),
            .I(N__36918));
    Span4Mux_h I__7541 (
            .O(N__36918),
            .I(N__36915));
    Odrv4 I__7540 (
            .O(N__36915),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__7539 (
            .O(N__36912),
            .I(N__36907));
    InMux I__7538 (
            .O(N__36911),
            .I(N__36902));
    InMux I__7537 (
            .O(N__36910),
            .I(N__36902));
    LocalMux I__7536 (
            .O(N__36907),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__7535 (
            .O(N__36902),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__7534 (
            .O(N__36897),
            .I(N__36894));
    InMux I__7533 (
            .O(N__36894),
            .I(N__36888));
    InMux I__7532 (
            .O(N__36893),
            .I(N__36888));
    LocalMux I__7531 (
            .O(N__36888),
            .I(N__36885));
    Odrv4 I__7530 (
            .O(N__36885),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__7529 (
            .O(N__36882),
            .I(N__36875));
    InMux I__7528 (
            .O(N__36881),
            .I(N__36875));
    InMux I__7527 (
            .O(N__36880),
            .I(N__36872));
    LocalMux I__7526 (
            .O(N__36875),
            .I(N__36869));
    LocalMux I__7525 (
            .O(N__36872),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__7524 (
            .O(N__36869),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__7523 (
            .O(N__36864),
            .I(N__36861));
    LocalMux I__7522 (
            .O(N__36861),
            .I(N__36858));
    Span4Mux_v I__7521 (
            .O(N__36858),
            .I(N__36855));
    Odrv4 I__7520 (
            .O(N__36855),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    CascadeMux I__7519 (
            .O(N__36852),
            .I(N__36849));
    InMux I__7518 (
            .O(N__36849),
            .I(N__36846));
    LocalMux I__7517 (
            .O(N__36846),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    CascadeMux I__7516 (
            .O(N__36843),
            .I(N__36840));
    InMux I__7515 (
            .O(N__36840),
            .I(N__36837));
    LocalMux I__7514 (
            .O(N__36837),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    CascadeMux I__7513 (
            .O(N__36834),
            .I(N__36831));
    InMux I__7512 (
            .O(N__36831),
            .I(N__36828));
    LocalMux I__7511 (
            .O(N__36828),
            .I(N__36825));
    Odrv4 I__7510 (
            .O(N__36825),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    InMux I__7509 (
            .O(N__36822),
            .I(N__36819));
    LocalMux I__7508 (
            .O(N__36819),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__7507 (
            .O(N__36816),
            .I(N__36813));
    LocalMux I__7506 (
            .O(N__36813),
            .I(N__36810));
    Odrv12 I__7505 (
            .O(N__36810),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__7504 (
            .O(N__36807),
            .I(N__36804));
    LocalMux I__7503 (
            .O(N__36804),
            .I(N__36801));
    Span4Mux_h I__7502 (
            .O(N__36801),
            .I(N__36798));
    Odrv4 I__7501 (
            .O(N__36798),
            .I(\current_shift_inst.control_input_axb_21 ));
    InMux I__7500 (
            .O(N__36795),
            .I(N__36791));
    InMux I__7499 (
            .O(N__36794),
            .I(N__36788));
    LocalMux I__7498 (
            .O(N__36791),
            .I(N__36785));
    LocalMux I__7497 (
            .O(N__36788),
            .I(N__36782));
    Span4Mux_h I__7496 (
            .O(N__36785),
            .I(N__36779));
    Odrv12 I__7495 (
            .O(N__36782),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    Odrv4 I__7494 (
            .O(N__36779),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__7493 (
            .O(N__36774),
            .I(N__36770));
    InMux I__7492 (
            .O(N__36773),
            .I(N__36767));
    LocalMux I__7491 (
            .O(N__36770),
            .I(N__36764));
    LocalMux I__7490 (
            .O(N__36767),
            .I(N__36759));
    Span4Mux_h I__7489 (
            .O(N__36764),
            .I(N__36756));
    InMux I__7488 (
            .O(N__36763),
            .I(N__36753));
    InMux I__7487 (
            .O(N__36762),
            .I(N__36750));
    Span4Mux_v I__7486 (
            .O(N__36759),
            .I(N__36747));
    Span4Mux_v I__7485 (
            .O(N__36756),
            .I(N__36744));
    LocalMux I__7484 (
            .O(N__36753),
            .I(N__36741));
    LocalMux I__7483 (
            .O(N__36750),
            .I(N__36738));
    Span4Mux_v I__7482 (
            .O(N__36747),
            .I(N__36733));
    Span4Mux_v I__7481 (
            .O(N__36744),
            .I(N__36733));
    Span4Mux_h I__7480 (
            .O(N__36741),
            .I(N__36728));
    Span4Mux_v I__7479 (
            .O(N__36738),
            .I(N__36728));
    Odrv4 I__7478 (
            .O(N__36733),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__7477 (
            .O(N__36728),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__7476 (
            .O(N__36723),
            .I(N__36715));
    CascadeMux I__7475 (
            .O(N__36722),
            .I(N__36708));
    CascadeMux I__7474 (
            .O(N__36721),
            .I(N__36705));
    InMux I__7473 (
            .O(N__36720),
            .I(N__36695));
    InMux I__7472 (
            .O(N__36719),
            .I(N__36695));
    InMux I__7471 (
            .O(N__36718),
            .I(N__36692));
    LocalMux I__7470 (
            .O(N__36715),
            .I(N__36683));
    InMux I__7469 (
            .O(N__36714),
            .I(N__36667));
    InMux I__7468 (
            .O(N__36713),
            .I(N__36664));
    InMux I__7467 (
            .O(N__36712),
            .I(N__36659));
    InMux I__7466 (
            .O(N__36711),
            .I(N__36659));
    InMux I__7465 (
            .O(N__36708),
            .I(N__36652));
    InMux I__7464 (
            .O(N__36705),
            .I(N__36652));
    InMux I__7463 (
            .O(N__36704),
            .I(N__36652));
    CascadeMux I__7462 (
            .O(N__36703),
            .I(N__36646));
    InMux I__7461 (
            .O(N__36702),
            .I(N__36642));
    InMux I__7460 (
            .O(N__36701),
            .I(N__36625));
    InMux I__7459 (
            .O(N__36700),
            .I(N__36625));
    LocalMux I__7458 (
            .O(N__36695),
            .I(N__36620));
    LocalMux I__7457 (
            .O(N__36692),
            .I(N__36620));
    InMux I__7456 (
            .O(N__36691),
            .I(N__36613));
    InMux I__7455 (
            .O(N__36690),
            .I(N__36613));
    InMux I__7454 (
            .O(N__36689),
            .I(N__36613));
    InMux I__7453 (
            .O(N__36688),
            .I(N__36610));
    InMux I__7452 (
            .O(N__36687),
            .I(N__36607));
    InMux I__7451 (
            .O(N__36686),
            .I(N__36604));
    Span4Mux_h I__7450 (
            .O(N__36683),
            .I(N__36599));
    InMux I__7449 (
            .O(N__36682),
            .I(N__36594));
    InMux I__7448 (
            .O(N__36681),
            .I(N__36591));
    InMux I__7447 (
            .O(N__36680),
            .I(N__36586));
    InMux I__7446 (
            .O(N__36679),
            .I(N__36586));
    InMux I__7445 (
            .O(N__36678),
            .I(N__36573));
    InMux I__7444 (
            .O(N__36677),
            .I(N__36573));
    InMux I__7443 (
            .O(N__36676),
            .I(N__36573));
    InMux I__7442 (
            .O(N__36675),
            .I(N__36573));
    InMux I__7441 (
            .O(N__36674),
            .I(N__36573));
    InMux I__7440 (
            .O(N__36673),
            .I(N__36573));
    InMux I__7439 (
            .O(N__36672),
            .I(N__36570));
    InMux I__7438 (
            .O(N__36671),
            .I(N__36565));
    InMux I__7437 (
            .O(N__36670),
            .I(N__36565));
    LocalMux I__7436 (
            .O(N__36667),
            .I(N__36562));
    LocalMux I__7435 (
            .O(N__36664),
            .I(N__36550));
    LocalMux I__7434 (
            .O(N__36659),
            .I(N__36550));
    LocalMux I__7433 (
            .O(N__36652),
            .I(N__36547));
    InMux I__7432 (
            .O(N__36651),
            .I(N__36539));
    InMux I__7431 (
            .O(N__36650),
            .I(N__36530));
    InMux I__7430 (
            .O(N__36649),
            .I(N__36530));
    InMux I__7429 (
            .O(N__36646),
            .I(N__36530));
    InMux I__7428 (
            .O(N__36645),
            .I(N__36530));
    LocalMux I__7427 (
            .O(N__36642),
            .I(N__36527));
    InMux I__7426 (
            .O(N__36641),
            .I(N__36518));
    InMux I__7425 (
            .O(N__36640),
            .I(N__36518));
    InMux I__7424 (
            .O(N__36639),
            .I(N__36518));
    InMux I__7423 (
            .O(N__36638),
            .I(N__36518));
    InMux I__7422 (
            .O(N__36637),
            .I(N__36513));
    InMux I__7421 (
            .O(N__36636),
            .I(N__36513));
    InMux I__7420 (
            .O(N__36635),
            .I(N__36506));
    InMux I__7419 (
            .O(N__36634),
            .I(N__36506));
    InMux I__7418 (
            .O(N__36633),
            .I(N__36506));
    InMux I__7417 (
            .O(N__36632),
            .I(N__36503));
    InMux I__7416 (
            .O(N__36631),
            .I(N__36498));
    InMux I__7415 (
            .O(N__36630),
            .I(N__36498));
    LocalMux I__7414 (
            .O(N__36625),
            .I(N__36491));
    Span4Mux_v I__7413 (
            .O(N__36620),
            .I(N__36491));
    LocalMux I__7412 (
            .O(N__36613),
            .I(N__36491));
    LocalMux I__7411 (
            .O(N__36610),
            .I(N__36484));
    LocalMux I__7410 (
            .O(N__36607),
            .I(N__36484));
    LocalMux I__7409 (
            .O(N__36604),
            .I(N__36484));
    InMux I__7408 (
            .O(N__36603),
            .I(N__36479));
    InMux I__7407 (
            .O(N__36602),
            .I(N__36479));
    Span4Mux_h I__7406 (
            .O(N__36599),
            .I(N__36474));
    InMux I__7405 (
            .O(N__36598),
            .I(N__36457));
    InMux I__7404 (
            .O(N__36597),
            .I(N__36457));
    LocalMux I__7403 (
            .O(N__36594),
            .I(N__36454));
    LocalMux I__7402 (
            .O(N__36591),
            .I(N__36451));
    LocalMux I__7401 (
            .O(N__36586),
            .I(N__36446));
    LocalMux I__7400 (
            .O(N__36573),
            .I(N__36446));
    LocalMux I__7399 (
            .O(N__36570),
            .I(N__36439));
    LocalMux I__7398 (
            .O(N__36565),
            .I(N__36439));
    Span4Mux_v I__7397 (
            .O(N__36562),
            .I(N__36439));
    InMux I__7396 (
            .O(N__36561),
            .I(N__36432));
    InMux I__7395 (
            .O(N__36560),
            .I(N__36432));
    InMux I__7394 (
            .O(N__36559),
            .I(N__36432));
    InMux I__7393 (
            .O(N__36558),
            .I(N__36423));
    InMux I__7392 (
            .O(N__36557),
            .I(N__36423));
    InMux I__7391 (
            .O(N__36556),
            .I(N__36423));
    InMux I__7390 (
            .O(N__36555),
            .I(N__36423));
    Span4Mux_h I__7389 (
            .O(N__36550),
            .I(N__36418));
    Span4Mux_s3_v I__7388 (
            .O(N__36547),
            .I(N__36418));
    InMux I__7387 (
            .O(N__36546),
            .I(N__36401));
    InMux I__7386 (
            .O(N__36545),
            .I(N__36401));
    InMux I__7385 (
            .O(N__36544),
            .I(N__36394));
    InMux I__7384 (
            .O(N__36543),
            .I(N__36394));
    InMux I__7383 (
            .O(N__36542),
            .I(N__36394));
    LocalMux I__7382 (
            .O(N__36539),
            .I(N__36391));
    LocalMux I__7381 (
            .O(N__36530),
            .I(N__36378));
    Span4Mux_h I__7380 (
            .O(N__36527),
            .I(N__36378));
    LocalMux I__7379 (
            .O(N__36518),
            .I(N__36378));
    LocalMux I__7378 (
            .O(N__36513),
            .I(N__36378));
    LocalMux I__7377 (
            .O(N__36506),
            .I(N__36378));
    LocalMux I__7376 (
            .O(N__36503),
            .I(N__36378));
    LocalMux I__7375 (
            .O(N__36498),
            .I(N__36371));
    Span4Mux_v I__7374 (
            .O(N__36491),
            .I(N__36371));
    Span4Mux_v I__7373 (
            .O(N__36484),
            .I(N__36371));
    LocalMux I__7372 (
            .O(N__36479),
            .I(N__36368));
    InMux I__7371 (
            .O(N__36478),
            .I(N__36365));
    InMux I__7370 (
            .O(N__36477),
            .I(N__36362));
    Span4Mux_v I__7369 (
            .O(N__36474),
            .I(N__36359));
    InMux I__7368 (
            .O(N__36473),
            .I(N__36356));
    InMux I__7367 (
            .O(N__36472),
            .I(N__36353));
    InMux I__7366 (
            .O(N__36471),
            .I(N__36346));
    InMux I__7365 (
            .O(N__36470),
            .I(N__36346));
    InMux I__7364 (
            .O(N__36469),
            .I(N__36346));
    InMux I__7363 (
            .O(N__36468),
            .I(N__36341));
    InMux I__7362 (
            .O(N__36467),
            .I(N__36341));
    InMux I__7361 (
            .O(N__36466),
            .I(N__36330));
    InMux I__7360 (
            .O(N__36465),
            .I(N__36330));
    InMux I__7359 (
            .O(N__36464),
            .I(N__36330));
    InMux I__7358 (
            .O(N__36463),
            .I(N__36330));
    InMux I__7357 (
            .O(N__36462),
            .I(N__36330));
    LocalMux I__7356 (
            .O(N__36457),
            .I(N__36327));
    Span4Mux_v I__7355 (
            .O(N__36454),
            .I(N__36318));
    Span4Mux_v I__7354 (
            .O(N__36451),
            .I(N__36318));
    Span4Mux_v I__7353 (
            .O(N__36446),
            .I(N__36318));
    Span4Mux_v I__7352 (
            .O(N__36439),
            .I(N__36318));
    LocalMux I__7351 (
            .O(N__36432),
            .I(N__36311));
    LocalMux I__7350 (
            .O(N__36423),
            .I(N__36311));
    Span4Mux_v I__7349 (
            .O(N__36418),
            .I(N__36311));
    InMux I__7348 (
            .O(N__36417),
            .I(N__36302));
    InMux I__7347 (
            .O(N__36416),
            .I(N__36302));
    InMux I__7346 (
            .O(N__36415),
            .I(N__36302));
    InMux I__7345 (
            .O(N__36414),
            .I(N__36302));
    InMux I__7344 (
            .O(N__36413),
            .I(N__36291));
    InMux I__7343 (
            .O(N__36412),
            .I(N__36291));
    InMux I__7342 (
            .O(N__36411),
            .I(N__36291));
    InMux I__7341 (
            .O(N__36410),
            .I(N__36291));
    InMux I__7340 (
            .O(N__36409),
            .I(N__36291));
    InMux I__7339 (
            .O(N__36408),
            .I(N__36284));
    InMux I__7338 (
            .O(N__36407),
            .I(N__36284));
    InMux I__7337 (
            .O(N__36406),
            .I(N__36284));
    LocalMux I__7336 (
            .O(N__36401),
            .I(N__36273));
    LocalMux I__7335 (
            .O(N__36394),
            .I(N__36273));
    Span4Mux_h I__7334 (
            .O(N__36391),
            .I(N__36273));
    Span4Mux_v I__7333 (
            .O(N__36378),
            .I(N__36273));
    Span4Mux_h I__7332 (
            .O(N__36371),
            .I(N__36273));
    Span4Mux_v I__7331 (
            .O(N__36368),
            .I(N__36264));
    LocalMux I__7330 (
            .O(N__36365),
            .I(N__36264));
    LocalMux I__7329 (
            .O(N__36362),
            .I(N__36264));
    Span4Mux_v I__7328 (
            .O(N__36359),
            .I(N__36264));
    LocalMux I__7327 (
            .O(N__36356),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__7326 (
            .O(N__36353),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__7325 (
            .O(N__36346),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__7324 (
            .O(N__36341),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__7323 (
            .O(N__36330),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__7322 (
            .O(N__36327),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__7321 (
            .O(N__36318),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__7320 (
            .O(N__36311),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__7319 (
            .O(N__36302),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__7318 (
            .O(N__36291),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__7317 (
            .O(N__36284),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__7316 (
            .O(N__36273),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__7315 (
            .O(N__36264),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__7314 (
            .O(N__36237),
            .I(N__36234));
    LocalMux I__7313 (
            .O(N__36234),
            .I(N__36231));
    Span4Mux_h I__7312 (
            .O(N__36231),
            .I(N__36227));
    InMux I__7311 (
            .O(N__36230),
            .I(N__36224));
    Span4Mux_v I__7310 (
            .O(N__36227),
            .I(N__36220));
    LocalMux I__7309 (
            .O(N__36224),
            .I(N__36217));
    InMux I__7308 (
            .O(N__36223),
            .I(N__36214));
    Sp12to4 I__7307 (
            .O(N__36220),
            .I(N__36209));
    Span12Mux_h I__7306 (
            .O(N__36217),
            .I(N__36209));
    LocalMux I__7305 (
            .O(N__36214),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    Odrv12 I__7304 (
            .O(N__36209),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    InMux I__7303 (
            .O(N__36204),
            .I(N__36201));
    LocalMux I__7302 (
            .O(N__36201),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__7301 (
            .O(N__36198),
            .I(N__36192));
    InMux I__7300 (
            .O(N__36197),
            .I(N__36189));
    InMux I__7299 (
            .O(N__36196),
            .I(N__36184));
    InMux I__7298 (
            .O(N__36195),
            .I(N__36184));
    LocalMux I__7297 (
            .O(N__36192),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7296 (
            .O(N__36189),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7295 (
            .O(N__36184),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__7294 (
            .O(N__36177),
            .I(N__36174));
    LocalMux I__7293 (
            .O(N__36174),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    CascadeMux I__7292 (
            .O(N__36171),
            .I(N__36168));
    InMux I__7291 (
            .O(N__36168),
            .I(N__36165));
    LocalMux I__7290 (
            .O(N__36165),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__7289 (
            .O(N__36162),
            .I(N__36159));
    LocalMux I__7288 (
            .O(N__36159),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    CascadeMux I__7287 (
            .O(N__36156),
            .I(N__36153));
    InMux I__7286 (
            .O(N__36153),
            .I(N__36150));
    LocalMux I__7285 (
            .O(N__36150),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__7284 (
            .O(N__36147),
            .I(N__36144));
    LocalMux I__7283 (
            .O(N__36144),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    CascadeMux I__7282 (
            .O(N__36141),
            .I(N__36138));
    InMux I__7281 (
            .O(N__36138),
            .I(N__36135));
    LocalMux I__7280 (
            .O(N__36135),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    InMux I__7279 (
            .O(N__36132),
            .I(N__36129));
    LocalMux I__7278 (
            .O(N__36129),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__7277 (
            .O(N__36126),
            .I(N__36123));
    LocalMux I__7276 (
            .O(N__36123),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__7275 (
            .O(N__36120),
            .I(N__36117));
    LocalMux I__7274 (
            .O(N__36117),
            .I(N__36114));
    Odrv4 I__7273 (
            .O(N__36114),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__7272 (
            .O(N__36111),
            .I(N__36108));
    LocalMux I__7271 (
            .O(N__36108),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__7270 (
            .O(N__36105),
            .I(N__36102));
    LocalMux I__7269 (
            .O(N__36102),
            .I(N__36099));
    Span4Mux_h I__7268 (
            .O(N__36099),
            .I(N__36096));
    Odrv4 I__7267 (
            .O(N__36096),
            .I(\current_shift_inst.control_input_axb_22 ));
    InMux I__7266 (
            .O(N__36093),
            .I(N__36090));
    LocalMux I__7265 (
            .O(N__36090),
            .I(N__36087));
    Span4Mux_v I__7264 (
            .O(N__36087),
            .I(N__36084));
    Odrv4 I__7263 (
            .O(N__36084),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__7262 (
            .O(N__36081),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__7261 (
            .O(N__36078),
            .I(N__36075));
    LocalMux I__7260 (
            .O(N__36075),
            .I(N__36072));
    Span4Mux_v I__7259 (
            .O(N__36072),
            .I(N__36069));
    Odrv4 I__7258 (
            .O(N__36069),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__7257 (
            .O(N__36066),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__7256 (
            .O(N__36063),
            .I(N__36060));
    LocalMux I__7255 (
            .O(N__36060),
            .I(N__36057));
    Span4Mux_h I__7254 (
            .O(N__36057),
            .I(N__36054));
    Odrv4 I__7253 (
            .O(N__36054),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__7252 (
            .O(N__36051),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__7251 (
            .O(N__36048),
            .I(N__36045));
    LocalMux I__7250 (
            .O(N__36045),
            .I(N__36042));
    Odrv4 I__7249 (
            .O(N__36042),
            .I(\current_shift_inst.control_input_axb_28 ));
    InMux I__7248 (
            .O(N__36039),
            .I(N__36036));
    LocalMux I__7247 (
            .O(N__36036),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    CascadeMux I__7246 (
            .O(N__36033),
            .I(N__36030));
    InMux I__7245 (
            .O(N__36030),
            .I(N__36027));
    LocalMux I__7244 (
            .O(N__36027),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    InMux I__7243 (
            .O(N__36024),
            .I(N__36021));
    LocalMux I__7242 (
            .O(N__36021),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    InMux I__7241 (
            .O(N__36018),
            .I(N__36015));
    LocalMux I__7240 (
            .O(N__36015),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__7239 (
            .O(N__36012),
            .I(N__36009));
    LocalMux I__7238 (
            .O(N__36009),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    InMux I__7237 (
            .O(N__36006),
            .I(N__36003));
    LocalMux I__7236 (
            .O(N__36003),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__7235 (
            .O(N__36000),
            .I(N__35997));
    LocalMux I__7234 (
            .O(N__35997),
            .I(N__35994));
    Span4Mux_v I__7233 (
            .O(N__35994),
            .I(N__35991));
    Odrv4 I__7232 (
            .O(N__35991),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__7231 (
            .O(N__35988),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__7230 (
            .O(N__35985),
            .I(N__35982));
    LocalMux I__7229 (
            .O(N__35982),
            .I(N__35979));
    Span4Mux_h I__7228 (
            .O(N__35979),
            .I(N__35976));
    Odrv4 I__7227 (
            .O(N__35976),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__7226 (
            .O(N__35973),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__7225 (
            .O(N__35970),
            .I(N__35967));
    LocalMux I__7224 (
            .O(N__35967),
            .I(N__35964));
    Span4Mux_h I__7223 (
            .O(N__35964),
            .I(N__35961));
    Odrv4 I__7222 (
            .O(N__35961),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__7221 (
            .O(N__35958),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__7220 (
            .O(N__35955),
            .I(bfn_14_16_0_));
    InMux I__7219 (
            .O(N__35952),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__7218 (
            .O(N__35949),
            .I(N__35946));
    LocalMux I__7217 (
            .O(N__35946),
            .I(N__35943));
    Odrv4 I__7216 (
            .O(N__35943),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__7215 (
            .O(N__35940),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__7214 (
            .O(N__35937),
            .I(N__35934));
    LocalMux I__7213 (
            .O(N__35934),
            .I(N__35931));
    Odrv4 I__7212 (
            .O(N__35931),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__7211 (
            .O(N__35928),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__7210 (
            .O(N__35925),
            .I(N__35922));
    LocalMux I__7209 (
            .O(N__35922),
            .I(N__35919));
    Span4Mux_v I__7208 (
            .O(N__35919),
            .I(N__35916));
    Odrv4 I__7207 (
            .O(N__35916),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__7206 (
            .O(N__35913),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__7205 (
            .O(N__35910),
            .I(N__35907));
    LocalMux I__7204 (
            .O(N__35907),
            .I(N__35904));
    Span4Mux_v I__7203 (
            .O(N__35904),
            .I(N__35901));
    Odrv4 I__7202 (
            .O(N__35901),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__7201 (
            .O(N__35898),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__7200 (
            .O(N__35895),
            .I(N__35892));
    LocalMux I__7199 (
            .O(N__35892),
            .I(N__35889));
    Span4Mux_h I__7198 (
            .O(N__35889),
            .I(N__35886));
    Odrv4 I__7197 (
            .O(N__35886),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__7196 (
            .O(N__35883),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    InMux I__7195 (
            .O(N__35880),
            .I(N__35877));
    LocalMux I__7194 (
            .O(N__35877),
            .I(N__35874));
    Span4Mux_h I__7193 (
            .O(N__35874),
            .I(N__35871));
    Odrv4 I__7192 (
            .O(N__35871),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__7191 (
            .O(N__35868),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__7190 (
            .O(N__35865),
            .I(N__35862));
    LocalMux I__7189 (
            .O(N__35862),
            .I(N__35859));
    Span4Mux_h I__7188 (
            .O(N__35859),
            .I(N__35856));
    Odrv4 I__7187 (
            .O(N__35856),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__7186 (
            .O(N__35853),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    InMux I__7185 (
            .O(N__35850),
            .I(N__35847));
    LocalMux I__7184 (
            .O(N__35847),
            .I(N__35844));
    Odrv4 I__7183 (
            .O(N__35844),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__7182 (
            .O(N__35841),
            .I(bfn_14_15_0_));
    InMux I__7181 (
            .O(N__35838),
            .I(N__35835));
    LocalMux I__7180 (
            .O(N__35835),
            .I(N__35832));
    Odrv4 I__7179 (
            .O(N__35832),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__7178 (
            .O(N__35829),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    InMux I__7177 (
            .O(N__35826),
            .I(N__35823));
    LocalMux I__7176 (
            .O(N__35823),
            .I(N__35820));
    Odrv4 I__7175 (
            .O(N__35820),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__7174 (
            .O(N__35817),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__7173 (
            .O(N__35814),
            .I(N__35811));
    LocalMux I__7172 (
            .O(N__35811),
            .I(N__35808));
    Span4Mux_h I__7171 (
            .O(N__35808),
            .I(N__35805));
    Odrv4 I__7170 (
            .O(N__35805),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__7169 (
            .O(N__35802),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    InMux I__7168 (
            .O(N__35799),
            .I(N__35796));
    LocalMux I__7167 (
            .O(N__35796),
            .I(N__35793));
    Span4Mux_h I__7166 (
            .O(N__35793),
            .I(N__35790));
    Odrv4 I__7165 (
            .O(N__35790),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__7164 (
            .O(N__35787),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__7163 (
            .O(N__35784),
            .I(\current_shift_inst.un38_control_input_cry_2_s0 ));
    InMux I__7162 (
            .O(N__35781),
            .I(\current_shift_inst.un38_control_input_cry_3_s0 ));
    InMux I__7161 (
            .O(N__35778),
            .I(N__35775));
    LocalMux I__7160 (
            .O(N__35775),
            .I(N__35772));
    Span4Mux_h I__7159 (
            .O(N__35772),
            .I(N__35769));
    Odrv4 I__7158 (
            .O(N__35769),
            .I(\current_shift_inst.un38_control_input_0_s0_5 ));
    InMux I__7157 (
            .O(N__35766),
            .I(\current_shift_inst.un38_control_input_cry_4_s0 ));
    InMux I__7156 (
            .O(N__35763),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__7155 (
            .O(N__35760),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    InMux I__7154 (
            .O(N__35757),
            .I(bfn_14_14_0_));
    InMux I__7153 (
            .O(N__35754),
            .I(N__35751));
    LocalMux I__7152 (
            .O(N__35751),
            .I(N__35748));
    Span4Mux_h I__7151 (
            .O(N__35748),
            .I(N__35745));
    Odrv4 I__7150 (
            .O(N__35745),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__7149 (
            .O(N__35742),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    InMux I__7148 (
            .O(N__35739),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__7147 (
            .O(N__35736),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    CascadeMux I__7146 (
            .O(N__35733),
            .I(N__35730));
    InMux I__7145 (
            .O(N__35730),
            .I(N__35727));
    LocalMux I__7144 (
            .O(N__35727),
            .I(N__35724));
    Span4Mux_v I__7143 (
            .O(N__35724),
            .I(N__35721));
    Odrv4 I__7142 (
            .O(N__35721),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    InMux I__7141 (
            .O(N__35718),
            .I(N__35714));
    InMux I__7140 (
            .O(N__35717),
            .I(N__35711));
    LocalMux I__7139 (
            .O(N__35714),
            .I(N__35707));
    LocalMux I__7138 (
            .O(N__35711),
            .I(N__35702));
    InMux I__7137 (
            .O(N__35710),
            .I(N__35699));
    Span4Mux_h I__7136 (
            .O(N__35707),
            .I(N__35696));
    InMux I__7135 (
            .O(N__35706),
            .I(N__35691));
    InMux I__7134 (
            .O(N__35705),
            .I(N__35691));
    Span4Mux_v I__7133 (
            .O(N__35702),
            .I(N__35688));
    LocalMux I__7132 (
            .O(N__35699),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__7131 (
            .O(N__35696),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__7130 (
            .O(N__35691),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__7129 (
            .O(N__35688),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__7128 (
            .O(N__35679),
            .I(N__35675));
    InMux I__7127 (
            .O(N__35678),
            .I(N__35672));
    LocalMux I__7126 (
            .O(N__35675),
            .I(N__35669));
    LocalMux I__7125 (
            .O(N__35672),
            .I(N__35664));
    Span4Mux_v I__7124 (
            .O(N__35669),
            .I(N__35664));
    Odrv4 I__7123 (
            .O(N__35664),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__7122 (
            .O(N__35661),
            .I(N__35657));
    InMux I__7121 (
            .O(N__35660),
            .I(N__35652));
    LocalMux I__7120 (
            .O(N__35657),
            .I(N__35649));
    CascadeMux I__7119 (
            .O(N__35656),
            .I(N__35646));
    InMux I__7118 (
            .O(N__35655),
            .I(N__35643));
    LocalMux I__7117 (
            .O(N__35652),
            .I(N__35638));
    Span4Mux_h I__7116 (
            .O(N__35649),
            .I(N__35638));
    InMux I__7115 (
            .O(N__35646),
            .I(N__35635));
    LocalMux I__7114 (
            .O(N__35643),
            .I(N__35632));
    Span4Mux_v I__7113 (
            .O(N__35638),
            .I(N__35629));
    LocalMux I__7112 (
            .O(N__35635),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__7111 (
            .O(N__35632),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__7110 (
            .O(N__35629),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__7109 (
            .O(N__35622),
            .I(N__35613));
    InMux I__7108 (
            .O(N__35621),
            .I(N__35613));
    InMux I__7107 (
            .O(N__35620),
            .I(N__35606));
    InMux I__7106 (
            .O(N__35619),
            .I(N__35606));
    InMux I__7105 (
            .O(N__35618),
            .I(N__35606));
    LocalMux I__7104 (
            .O(N__35613),
            .I(N__35603));
    LocalMux I__7103 (
            .O(N__35606),
            .I(N__35600));
    Span12Mux_s11_v I__7102 (
            .O(N__35603),
            .I(N__35597));
    Span4Mux_h I__7101 (
            .O(N__35600),
            .I(N__35594));
    Odrv12 I__7100 (
            .O(N__35597),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__7099 (
            .O(N__35594),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__7098 (
            .O(N__35589),
            .I(N__35586));
    LocalMux I__7097 (
            .O(N__35586),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    CascadeMux I__7096 (
            .O(N__35583),
            .I(N__35578));
    InMux I__7095 (
            .O(N__35582),
            .I(N__35575));
    InMux I__7094 (
            .O(N__35581),
            .I(N__35570));
    InMux I__7093 (
            .O(N__35578),
            .I(N__35570));
    LocalMux I__7092 (
            .O(N__35575),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__7091 (
            .O(N__35570),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__7090 (
            .O(N__35565),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__7089 (
            .O(N__35562),
            .I(N__35555));
    InMux I__7088 (
            .O(N__35561),
            .I(N__35555));
    InMux I__7087 (
            .O(N__35560),
            .I(N__35552));
    LocalMux I__7086 (
            .O(N__35555),
            .I(N__35549));
    LocalMux I__7085 (
            .O(N__35552),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__7084 (
            .O(N__35549),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__7083 (
            .O(N__35544),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__7082 (
            .O(N__35541),
            .I(N__35534));
    InMux I__7081 (
            .O(N__35540),
            .I(N__35534));
    InMux I__7080 (
            .O(N__35539),
            .I(N__35531));
    LocalMux I__7079 (
            .O(N__35534),
            .I(N__35528));
    LocalMux I__7078 (
            .O(N__35531),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__7077 (
            .O(N__35528),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__7076 (
            .O(N__35523),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    CascadeMux I__7075 (
            .O(N__35520),
            .I(N__35516));
    CascadeMux I__7074 (
            .O(N__35519),
            .I(N__35513));
    InMux I__7073 (
            .O(N__35516),
            .I(N__35510));
    InMux I__7072 (
            .O(N__35513),
            .I(N__35507));
    LocalMux I__7071 (
            .O(N__35510),
            .I(N__35503));
    LocalMux I__7070 (
            .O(N__35507),
            .I(N__35500));
    InMux I__7069 (
            .O(N__35506),
            .I(N__35497));
    Span4Mux_v I__7068 (
            .O(N__35503),
            .I(N__35494));
    Span4Mux_v I__7067 (
            .O(N__35500),
            .I(N__35491));
    LocalMux I__7066 (
            .O(N__35497),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__7065 (
            .O(N__35494),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__7064 (
            .O(N__35491),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__7063 (
            .O(N__35484),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__7062 (
            .O(N__35481),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__7061 (
            .O(N__35478),
            .I(N__35474));
    InMux I__7060 (
            .O(N__35477),
            .I(N__35471));
    LocalMux I__7059 (
            .O(N__35474),
            .I(N__35467));
    LocalMux I__7058 (
            .O(N__35471),
            .I(N__35464));
    InMux I__7057 (
            .O(N__35470),
            .I(N__35461));
    Span4Mux_v I__7056 (
            .O(N__35467),
            .I(N__35458));
    Span4Mux_v I__7055 (
            .O(N__35464),
            .I(N__35455));
    LocalMux I__7054 (
            .O(N__35461),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__7053 (
            .O(N__35458),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__7052 (
            .O(N__35455),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__7051 (
            .O(N__35448),
            .I(N__35445));
    LocalMux I__7050 (
            .O(N__35445),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    CascadeMux I__7049 (
            .O(N__35442),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ));
    InMux I__7048 (
            .O(N__35439),
            .I(N__35436));
    LocalMux I__7047 (
            .O(N__35436),
            .I(N__35433));
    Span4Mux_v I__7046 (
            .O(N__35433),
            .I(N__35430));
    Span4Mux_h I__7045 (
            .O(N__35430),
            .I(N__35427));
    Odrv4 I__7044 (
            .O(N__35427),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    CascadeMux I__7043 (
            .O(N__35424),
            .I(N__35421));
    InMux I__7042 (
            .O(N__35421),
            .I(N__35418));
    LocalMux I__7041 (
            .O(N__35418),
            .I(N__35415));
    Odrv4 I__7040 (
            .O(N__35415),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__7039 (
            .O(N__35412),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__7038 (
            .O(N__35409),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__7037 (
            .O(N__35406),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__7036 (
            .O(N__35403),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__7035 (
            .O(N__35400),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__7034 (
            .O(N__35397),
            .I(N__35390));
    InMux I__7033 (
            .O(N__35396),
            .I(N__35390));
    InMux I__7032 (
            .O(N__35395),
            .I(N__35387));
    LocalMux I__7031 (
            .O(N__35390),
            .I(N__35384));
    LocalMux I__7030 (
            .O(N__35387),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv12 I__7029 (
            .O(N__35384),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__7028 (
            .O(N__35379),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    CascadeMux I__7027 (
            .O(N__35376),
            .I(N__35372));
    InMux I__7026 (
            .O(N__35375),
            .I(N__35366));
    InMux I__7025 (
            .O(N__35372),
            .I(N__35366));
    InMux I__7024 (
            .O(N__35371),
            .I(N__35363));
    LocalMux I__7023 (
            .O(N__35366),
            .I(N__35360));
    LocalMux I__7022 (
            .O(N__35363),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv12 I__7021 (
            .O(N__35360),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__7020 (
            .O(N__35355),
            .I(bfn_14_10_0_));
    InMux I__7019 (
            .O(N__35352),
            .I(N__35347));
    InMux I__7018 (
            .O(N__35351),
            .I(N__35342));
    InMux I__7017 (
            .O(N__35350),
            .I(N__35342));
    LocalMux I__7016 (
            .O(N__35347),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__7015 (
            .O(N__35342),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__7014 (
            .O(N__35337),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__7013 (
            .O(N__35334),
            .I(N__35330));
    InMux I__7012 (
            .O(N__35333),
            .I(N__35327));
    LocalMux I__7011 (
            .O(N__35330),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__7010 (
            .O(N__35327),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__7009 (
            .O(N__35322),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__7008 (
            .O(N__35319),
            .I(N__35315));
    InMux I__7007 (
            .O(N__35318),
            .I(N__35312));
    LocalMux I__7006 (
            .O(N__35315),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__7005 (
            .O(N__35312),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__7004 (
            .O(N__35307),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__7003 (
            .O(N__35304),
            .I(N__35300));
    InMux I__7002 (
            .O(N__35303),
            .I(N__35297));
    LocalMux I__7001 (
            .O(N__35300),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__7000 (
            .O(N__35297),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__6999 (
            .O(N__35292),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__6998 (
            .O(N__35289),
            .I(N__35285));
    InMux I__6997 (
            .O(N__35288),
            .I(N__35282));
    LocalMux I__6996 (
            .O(N__35285),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__6995 (
            .O(N__35282),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__6994 (
            .O(N__35277),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__6993 (
            .O(N__35274),
            .I(N__35270));
    InMux I__6992 (
            .O(N__35273),
            .I(N__35267));
    LocalMux I__6991 (
            .O(N__35270),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__6990 (
            .O(N__35267),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__6989 (
            .O(N__35262),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__6988 (
            .O(N__35259),
            .I(N__35255));
    InMux I__6987 (
            .O(N__35258),
            .I(N__35252));
    LocalMux I__6986 (
            .O(N__35255),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__6985 (
            .O(N__35252),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__6984 (
            .O(N__35247),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__6983 (
            .O(N__35244),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__6982 (
            .O(N__35241),
            .I(bfn_14_9_0_));
    InMux I__6981 (
            .O(N__35238),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__6980 (
            .O(N__35235),
            .I(N__35231));
    InMux I__6979 (
            .O(N__35234),
            .I(N__35228));
    LocalMux I__6978 (
            .O(N__35231),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__6977 (
            .O(N__35228),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__6976 (
            .O(N__35223),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__6975 (
            .O(N__35220),
            .I(N__35217));
    InMux I__6974 (
            .O(N__35217),
            .I(N__35214));
    LocalMux I__6973 (
            .O(N__35214),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ));
    InMux I__6972 (
            .O(N__35211),
            .I(N__35207));
    InMux I__6971 (
            .O(N__35210),
            .I(N__35204));
    LocalMux I__6970 (
            .O(N__35207),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__6969 (
            .O(N__35204),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__6968 (
            .O(N__35199),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__6967 (
            .O(N__35196),
            .I(N__35192));
    InMux I__6966 (
            .O(N__35195),
            .I(N__35189));
    LocalMux I__6965 (
            .O(N__35192),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__6964 (
            .O(N__35189),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__6963 (
            .O(N__35184),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__6962 (
            .O(N__35181),
            .I(N__35177));
    InMux I__6961 (
            .O(N__35180),
            .I(N__35174));
    LocalMux I__6960 (
            .O(N__35177),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__6959 (
            .O(N__35174),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__6958 (
            .O(N__35169),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__6957 (
            .O(N__35166),
            .I(N__35162));
    InMux I__6956 (
            .O(N__35165),
            .I(N__35159));
    LocalMux I__6955 (
            .O(N__35162),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__6954 (
            .O(N__35159),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__6953 (
            .O(N__35154),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__6952 (
            .O(N__35151),
            .I(N__35147));
    InMux I__6951 (
            .O(N__35150),
            .I(N__35144));
    LocalMux I__6950 (
            .O(N__35147),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__6949 (
            .O(N__35144),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__6948 (
            .O(N__35139),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__6947 (
            .O(N__35136),
            .I(N__35132));
    InMux I__6946 (
            .O(N__35135),
            .I(N__35129));
    LocalMux I__6945 (
            .O(N__35132),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__6944 (
            .O(N__35129),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__6943 (
            .O(N__35124),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__6942 (
            .O(N__35121),
            .I(N__35117));
    InMux I__6941 (
            .O(N__35120),
            .I(N__35114));
    LocalMux I__6940 (
            .O(N__35117),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__6939 (
            .O(N__35114),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__6938 (
            .O(N__35109),
            .I(bfn_14_8_0_));
    InMux I__6937 (
            .O(N__35106),
            .I(N__35102));
    InMux I__6936 (
            .O(N__35105),
            .I(N__35099));
    LocalMux I__6935 (
            .O(N__35102),
            .I(N__35094));
    LocalMux I__6934 (
            .O(N__35099),
            .I(N__35094));
    Span4Mux_s3_v I__6933 (
            .O(N__35094),
            .I(N__35091));
    Span4Mux_h I__6932 (
            .O(N__35091),
            .I(N__35088));
    Sp12to4 I__6931 (
            .O(N__35088),
            .I(N__35079));
    InMux I__6930 (
            .O(N__35087),
            .I(N__35076));
    InMux I__6929 (
            .O(N__35086),
            .I(N__35071));
    InMux I__6928 (
            .O(N__35085),
            .I(N__35071));
    InMux I__6927 (
            .O(N__35084),
            .I(N__35064));
    InMux I__6926 (
            .O(N__35083),
            .I(N__35064));
    InMux I__6925 (
            .O(N__35082),
            .I(N__35064));
    Span12Mux_v I__6924 (
            .O(N__35079),
            .I(N__35061));
    LocalMux I__6923 (
            .O(N__35076),
            .I(N__35054));
    LocalMux I__6922 (
            .O(N__35071),
            .I(N__35054));
    LocalMux I__6921 (
            .O(N__35064),
            .I(N__35054));
    Span12Mux_v I__6920 (
            .O(N__35061),
            .I(N__35051));
    Span4Mux_v I__6919 (
            .O(N__35054),
            .I(N__35048));
    Span12Mux_h I__6918 (
            .O(N__35051),
            .I(N__35045));
    Span4Mux_h I__6917 (
            .O(N__35048),
            .I(N__35042));
    Odrv12 I__6916 (
            .O(N__35045),
            .I(start_stop_c));
    Odrv4 I__6915 (
            .O(N__35042),
            .I(start_stop_c));
    InMux I__6914 (
            .O(N__35037),
            .I(N__35032));
    InMux I__6913 (
            .O(N__35036),
            .I(N__35027));
    InMux I__6912 (
            .O(N__35035),
            .I(N__35027));
    LocalMux I__6911 (
            .O(N__35032),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    LocalMux I__6910 (
            .O(N__35027),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    CascadeMux I__6909 (
            .O(N__35022),
            .I(N__35018));
    InMux I__6908 (
            .O(N__35021),
            .I(N__35014));
    InMux I__6907 (
            .O(N__35018),
            .I(N__35009));
    InMux I__6906 (
            .O(N__35017),
            .I(N__35009));
    LocalMux I__6905 (
            .O(N__35014),
            .I(\phase_controller_inst2.start_flagZ0 ));
    LocalMux I__6904 (
            .O(N__35009),
            .I(\phase_controller_inst2.start_flagZ0 ));
    CascadeMux I__6903 (
            .O(N__35004),
            .I(N__35001));
    InMux I__6902 (
            .O(N__35001),
            .I(N__34998));
    LocalMux I__6901 (
            .O(N__34998),
            .I(N__34995));
    Span4Mux_v I__6900 (
            .O(N__34995),
            .I(N__34992));
    Odrv4 I__6899 (
            .O(N__34992),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    InMux I__6898 (
            .O(N__34989),
            .I(N__34986));
    LocalMux I__6897 (
            .O(N__34986),
            .I(N__34983));
    Span4Mux_v I__6896 (
            .O(N__34983),
            .I(N__34980));
    Odrv4 I__6895 (
            .O(N__34980),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    CascadeMux I__6894 (
            .O(N__34977),
            .I(elapsed_time_ns_1_RNIH33T9_0_5_cascade_));
    InMux I__6893 (
            .O(N__34974),
            .I(N__34971));
    LocalMux I__6892 (
            .O(N__34971),
            .I(N__34968));
    Odrv4 I__6891 (
            .O(N__34968),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__6890 (
            .O(N__34965),
            .I(elapsed_time_ns_1_RNI25DN9_0_24_cascade_));
    InMux I__6889 (
            .O(N__34962),
            .I(N__34956));
    InMux I__6888 (
            .O(N__34961),
            .I(N__34956));
    LocalMux I__6887 (
            .O(N__34956),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    InMux I__6886 (
            .O(N__34953),
            .I(N__34950));
    LocalMux I__6885 (
            .O(N__34950),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    CascadeMux I__6884 (
            .O(N__34947),
            .I(N__34943));
    InMux I__6883 (
            .O(N__34946),
            .I(N__34939));
    InMux I__6882 (
            .O(N__34943),
            .I(N__34936));
    InMux I__6881 (
            .O(N__34942),
            .I(N__34933));
    LocalMux I__6880 (
            .O(N__34939),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__6879 (
            .O(N__34936),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__6878 (
            .O(N__34933),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    IoInMux I__6877 (
            .O(N__34926),
            .I(N__34923));
    LocalMux I__6876 (
            .O(N__34923),
            .I(N__34920));
    Odrv12 I__6875 (
            .O(N__34920),
            .I(s2_phy_c));
    CascadeMux I__6874 (
            .O(N__34917),
            .I(N__34911));
    CascadeMux I__6873 (
            .O(N__34916),
            .I(N__34907));
    InMux I__6872 (
            .O(N__34915),
            .I(N__34902));
    InMux I__6871 (
            .O(N__34914),
            .I(N__34902));
    InMux I__6870 (
            .O(N__34911),
            .I(N__34899));
    CascadeMux I__6869 (
            .O(N__34910),
            .I(N__34896));
    InMux I__6868 (
            .O(N__34907),
            .I(N__34893));
    LocalMux I__6867 (
            .O(N__34902),
            .I(N__34888));
    LocalMux I__6866 (
            .O(N__34899),
            .I(N__34888));
    InMux I__6865 (
            .O(N__34896),
            .I(N__34884));
    LocalMux I__6864 (
            .O(N__34893),
            .I(N__34879));
    Span12Mux_v I__6863 (
            .O(N__34888),
            .I(N__34879));
    InMux I__6862 (
            .O(N__34887),
            .I(N__34876));
    LocalMux I__6861 (
            .O(N__34884),
            .I(state_3));
    Odrv12 I__6860 (
            .O(N__34879),
            .I(state_3));
    LocalMux I__6859 (
            .O(N__34876),
            .I(state_3));
    IoInMux I__6858 (
            .O(N__34869),
            .I(N__34866));
    LocalMux I__6857 (
            .O(N__34866),
            .I(N__34863));
    Span4Mux_s0_v I__6856 (
            .O(N__34863),
            .I(N__34860));
    Span4Mux_v I__6855 (
            .O(N__34860),
            .I(N__34857));
    Span4Mux_v I__6854 (
            .O(N__34857),
            .I(N__34852));
    InMux I__6853 (
            .O(N__34856),
            .I(N__34849));
    InMux I__6852 (
            .O(N__34855),
            .I(N__34846));
    Odrv4 I__6851 (
            .O(N__34852),
            .I(s1_phy_c));
    LocalMux I__6850 (
            .O(N__34849),
            .I(s1_phy_c));
    LocalMux I__6849 (
            .O(N__34846),
            .I(s1_phy_c));
    InMux I__6848 (
            .O(N__34839),
            .I(N__34833));
    InMux I__6847 (
            .O(N__34838),
            .I(N__34828));
    InMux I__6846 (
            .O(N__34837),
            .I(N__34828));
    InMux I__6845 (
            .O(N__34836),
            .I(N__34825));
    LocalMux I__6844 (
            .O(N__34833),
            .I(N__34822));
    LocalMux I__6843 (
            .O(N__34828),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6842 (
            .O(N__34825),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__6841 (
            .O(N__34822),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__6840 (
            .O(N__34815),
            .I(N__34807));
    InMux I__6839 (
            .O(N__34814),
            .I(N__34807));
    InMux I__6838 (
            .O(N__34813),
            .I(N__34804));
    InMux I__6837 (
            .O(N__34812),
            .I(N__34801));
    LocalMux I__6836 (
            .O(N__34807),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6835 (
            .O(N__34804),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6834 (
            .O(N__34801),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__6833 (
            .O(N__34794),
            .I(N__34791));
    LocalMux I__6832 (
            .O(N__34791),
            .I(N__34788));
    Span4Mux_s3_v I__6831 (
            .O(N__34788),
            .I(N__34785));
    Odrv4 I__6830 (
            .O(N__34785),
            .I(\current_shift_inst.timer_s1.N_161_i ));
    InMux I__6829 (
            .O(N__34782),
            .I(N__34779));
    LocalMux I__6828 (
            .O(N__34779),
            .I(N__34774));
    InMux I__6827 (
            .O(N__34778),
            .I(N__34771));
    InMux I__6826 (
            .O(N__34777),
            .I(N__34768));
    IoSpan4Mux I__6825 (
            .O(N__34774),
            .I(N__34765));
    LocalMux I__6824 (
            .O(N__34771),
            .I(N__34762));
    LocalMux I__6823 (
            .O(N__34768),
            .I(N__34759));
    IoSpan4Mux I__6822 (
            .O(N__34765),
            .I(N__34756));
    IoSpan4Mux I__6821 (
            .O(N__34762),
            .I(N__34751));
    IoSpan4Mux I__6820 (
            .O(N__34759),
            .I(N__34751));
    Odrv4 I__6819 (
            .O(N__34756),
            .I(il_min_comp1_c));
    Odrv4 I__6818 (
            .O(N__34751),
            .I(il_min_comp1_c));
    InMux I__6817 (
            .O(N__34746),
            .I(N__34742));
    InMux I__6816 (
            .O(N__34745),
            .I(N__34739));
    LocalMux I__6815 (
            .O(N__34742),
            .I(\phase_controller_inst1.N_61 ));
    LocalMux I__6814 (
            .O(N__34739),
            .I(\phase_controller_inst1.N_61 ));
    InMux I__6813 (
            .O(N__34734),
            .I(N__34731));
    LocalMux I__6812 (
            .O(N__34731),
            .I(N__34728));
    Sp12to4 I__6811 (
            .O(N__34728),
            .I(N__34723));
    InMux I__6810 (
            .O(N__34727),
            .I(N__34719));
    InMux I__6809 (
            .O(N__34726),
            .I(N__34716));
    Span12Mux_v I__6808 (
            .O(N__34723),
            .I(N__34713));
    InMux I__6807 (
            .O(N__34722),
            .I(N__34710));
    LocalMux I__6806 (
            .O(N__34719),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__6805 (
            .O(N__34716),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__6804 (
            .O(N__34713),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__6803 (
            .O(N__34710),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    InMux I__6802 (
            .O(N__34701),
            .I(bfn_13_19_0_));
    InMux I__6801 (
            .O(N__34698),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__6800 (
            .O(N__34695),
            .I(N__34692));
    LocalMux I__6799 (
            .O(N__34692),
            .I(N__34689));
    Odrv4 I__6798 (
            .O(N__34689),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__6797 (
            .O(N__34686),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__6796 (
            .O(N__34683),
            .I(N__34680));
    LocalMux I__6795 (
            .O(N__34680),
            .I(N__34677));
    Odrv4 I__6794 (
            .O(N__34677),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__6793 (
            .O(N__34674),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__6792 (
            .O(N__34671),
            .I(N__34668));
    LocalMux I__6791 (
            .O(N__34668),
            .I(N__34665));
    Odrv4 I__6790 (
            .O(N__34665),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__6789 (
            .O(N__34662),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__6788 (
            .O(N__34659),
            .I(N__34656));
    LocalMux I__6787 (
            .O(N__34656),
            .I(N__34653));
    Span4Mux_h I__6786 (
            .O(N__34653),
            .I(N__34650));
    Odrv4 I__6785 (
            .O(N__34650),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__6784 (
            .O(N__34647),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__6783 (
            .O(N__34644),
            .I(N__34641));
    LocalMux I__6782 (
            .O(N__34641),
            .I(N__34638));
    Span4Mux_h I__6781 (
            .O(N__34638),
            .I(N__34635));
    Odrv4 I__6780 (
            .O(N__34635),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__6779 (
            .O(N__34632),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__6778 (
            .O(N__34629),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__6777 (
            .O(N__34626),
            .I(N__34623));
    LocalMux I__6776 (
            .O(N__34623),
            .I(N__34620));
    Odrv4 I__6775 (
            .O(N__34620),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__6774 (
            .O(N__34617),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__6773 (
            .O(N__34614),
            .I(N__34611));
    LocalMux I__6772 (
            .O(N__34611),
            .I(N__34608));
    Odrv4 I__6771 (
            .O(N__34608),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    InMux I__6770 (
            .O(N__34605),
            .I(bfn_13_18_0_));
    InMux I__6769 (
            .O(N__34602),
            .I(N__34599));
    LocalMux I__6768 (
            .O(N__34599),
            .I(N__34596));
    Odrv4 I__6767 (
            .O(N__34596),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__6766 (
            .O(N__34593),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    InMux I__6765 (
            .O(N__34590),
            .I(N__34587));
    LocalMux I__6764 (
            .O(N__34587),
            .I(N__34584));
    Odrv4 I__6763 (
            .O(N__34584),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__6762 (
            .O(N__34581),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    InMux I__6761 (
            .O(N__34578),
            .I(N__34575));
    LocalMux I__6760 (
            .O(N__34575),
            .I(N__34572));
    Odrv4 I__6759 (
            .O(N__34572),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__6758 (
            .O(N__34569),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    InMux I__6757 (
            .O(N__34566),
            .I(N__34563));
    LocalMux I__6756 (
            .O(N__34563),
            .I(N__34560));
    Odrv4 I__6755 (
            .O(N__34560),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__6754 (
            .O(N__34557),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__6753 (
            .O(N__34554),
            .I(N__34551));
    LocalMux I__6752 (
            .O(N__34551),
            .I(N__34548));
    Odrv4 I__6751 (
            .O(N__34548),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__6750 (
            .O(N__34545),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__6749 (
            .O(N__34542),
            .I(N__34539));
    LocalMux I__6748 (
            .O(N__34539),
            .I(N__34536));
    Odrv4 I__6747 (
            .O(N__34536),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__6746 (
            .O(N__34533),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__6745 (
            .O(N__34530),
            .I(N__34527));
    LocalMux I__6744 (
            .O(N__34527),
            .I(N__34524));
    Odrv4 I__6743 (
            .O(N__34524),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__6742 (
            .O(N__34521),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__6741 (
            .O(N__34518),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    InMux I__6740 (
            .O(N__34515),
            .I(bfn_13_17_0_));
    InMux I__6739 (
            .O(N__34512),
            .I(N__34509));
    LocalMux I__6738 (
            .O(N__34509),
            .I(N__34506));
    Span4Mux_v I__6737 (
            .O(N__34506),
            .I(N__34503));
    Odrv4 I__6736 (
            .O(N__34503),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__6735 (
            .O(N__34500),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__6734 (
            .O(N__34497),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__6733 (
            .O(N__34494),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    InMux I__6732 (
            .O(N__34491),
            .I(N__34488));
    LocalMux I__6731 (
            .O(N__34488),
            .I(N__34485));
    Odrv4 I__6730 (
            .O(N__34485),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__6729 (
            .O(N__34482),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__6728 (
            .O(N__34479),
            .I(N__34476));
    LocalMux I__6727 (
            .O(N__34476),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__6726 (
            .O(N__34473),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    InMux I__6725 (
            .O(N__34470),
            .I(N__34467));
    LocalMux I__6724 (
            .O(N__34467),
            .I(N__34464));
    Odrv4 I__6723 (
            .O(N__34464),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__6722 (
            .O(N__34461),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    CascadeMux I__6721 (
            .O(N__34458),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    InMux I__6720 (
            .O(N__34455),
            .I(N__34450));
    InMux I__6719 (
            .O(N__34454),
            .I(N__34447));
    InMux I__6718 (
            .O(N__34453),
            .I(N__34444));
    LocalMux I__6717 (
            .O(N__34450),
            .I(N__34439));
    LocalMux I__6716 (
            .O(N__34447),
            .I(N__34439));
    LocalMux I__6715 (
            .O(N__34444),
            .I(N__34436));
    Odrv4 I__6714 (
            .O(N__34439),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__6713 (
            .O(N__34436),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__6712 (
            .O(N__34431),
            .I(N__34427));
    InMux I__6711 (
            .O(N__34430),
            .I(N__34424));
    LocalMux I__6710 (
            .O(N__34427),
            .I(N__34421));
    LocalMux I__6709 (
            .O(N__34424),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    Odrv4 I__6708 (
            .O(N__34421),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    InMux I__6707 (
            .O(N__34416),
            .I(N__34412));
    InMux I__6706 (
            .O(N__34415),
            .I(N__34409));
    LocalMux I__6705 (
            .O(N__34412),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    LocalMux I__6704 (
            .O(N__34409),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    CascadeMux I__6703 (
            .O(N__34404),
            .I(N__34401));
    InMux I__6702 (
            .O(N__34401),
            .I(N__34398));
    LocalMux I__6701 (
            .O(N__34398),
            .I(N__34395));
    Span4Mux_v I__6700 (
            .O(N__34395),
            .I(N__34392));
    Odrv4 I__6699 (
            .O(N__34392),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    InMux I__6698 (
            .O(N__34389),
            .I(\current_shift_inst.un38_control_input_cry_2_s1 ));
    InMux I__6697 (
            .O(N__34386),
            .I(\current_shift_inst.un38_control_input_cry_3_s1 ));
    InMux I__6696 (
            .O(N__34383),
            .I(N__34380));
    LocalMux I__6695 (
            .O(N__34380),
            .I(N__34377));
    Span4Mux_h I__6694 (
            .O(N__34377),
            .I(N__34374));
    Odrv4 I__6693 (
            .O(N__34374),
            .I(\current_shift_inst.un38_control_input_0_s1_5 ));
    InMux I__6692 (
            .O(N__34371),
            .I(\current_shift_inst.un38_control_input_cry_4_s1 ));
    InMux I__6691 (
            .O(N__34368),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__6690 (
            .O(N__34365),
            .I(N__34362));
    LocalMux I__6689 (
            .O(N__34362),
            .I(N__34359));
    Odrv12 I__6688 (
            .O(N__34359),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__6687 (
            .O(N__34356),
            .I(N__34353));
    LocalMux I__6686 (
            .O(N__34353),
            .I(N__34350));
    Odrv12 I__6685 (
            .O(N__34350),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__6684 (
            .O(N__34347),
            .I(N__34342));
    InMux I__6683 (
            .O(N__34346),
            .I(N__34339));
    InMux I__6682 (
            .O(N__34345),
            .I(N__34336));
    LocalMux I__6681 (
            .O(N__34342),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    LocalMux I__6680 (
            .O(N__34339),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    LocalMux I__6679 (
            .O(N__34336),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    InMux I__6678 (
            .O(N__34329),
            .I(N__34326));
    LocalMux I__6677 (
            .O(N__34326),
            .I(N__34323));
    Odrv12 I__6676 (
            .O(N__34323),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__6675 (
            .O(N__34320),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ));
    InMux I__6674 (
            .O(N__34317),
            .I(N__34314));
    LocalMux I__6673 (
            .O(N__34314),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    CascadeMux I__6672 (
            .O(N__34311),
            .I(N__34308));
    InMux I__6671 (
            .O(N__34308),
            .I(N__34305));
    LocalMux I__6670 (
            .O(N__34305),
            .I(N__34302));
    Odrv12 I__6669 (
            .O(N__34302),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__6668 (
            .O(N__34299),
            .I(N__34296));
    LocalMux I__6667 (
            .O(N__34296),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    CascadeMux I__6666 (
            .O(N__34293),
            .I(elapsed_time_ns_1_RNI47DN9_0_26_cascade_));
    InMux I__6665 (
            .O(N__34290),
            .I(N__34284));
    InMux I__6664 (
            .O(N__34289),
            .I(N__34284));
    LocalMux I__6663 (
            .O(N__34284),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    CascadeMux I__6662 (
            .O(N__34281),
            .I(N__34278));
    InMux I__6661 (
            .O(N__34278),
            .I(N__34275));
    LocalMux I__6660 (
            .O(N__34275),
            .I(N__34272));
    Odrv4 I__6659 (
            .O(N__34272),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__6658 (
            .O(N__34269),
            .I(N__34266));
    LocalMux I__6657 (
            .O(N__34266),
            .I(N__34262));
    InMux I__6656 (
            .O(N__34265),
            .I(N__34259));
    Odrv4 I__6655 (
            .O(N__34262),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__6654 (
            .O(N__34259),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    CascadeMux I__6653 (
            .O(N__34254),
            .I(elapsed_time_ns_1_RNI69DN9_0_28_cascade_));
    InMux I__6652 (
            .O(N__34251),
            .I(N__34247));
    InMux I__6651 (
            .O(N__34250),
            .I(N__34243));
    LocalMux I__6650 (
            .O(N__34247),
            .I(N__34240));
    InMux I__6649 (
            .O(N__34246),
            .I(N__34237));
    LocalMux I__6648 (
            .O(N__34243),
            .I(N__34234));
    Span4Mux_h I__6647 (
            .O(N__34240),
            .I(N__34231));
    LocalMux I__6646 (
            .O(N__34237),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    Odrv12 I__6645 (
            .O(N__34234),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    Odrv4 I__6644 (
            .O(N__34231),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    CascadeMux I__6643 (
            .O(N__34224),
            .I(N__34220));
    CascadeMux I__6642 (
            .O(N__34223),
            .I(N__34217));
    InMux I__6641 (
            .O(N__34220),
            .I(N__34212));
    InMux I__6640 (
            .O(N__34217),
            .I(N__34212));
    LocalMux I__6639 (
            .O(N__34212),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    InMux I__6638 (
            .O(N__34209),
            .I(N__34203));
    InMux I__6637 (
            .O(N__34208),
            .I(N__34203));
    LocalMux I__6636 (
            .O(N__34203),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    InMux I__6635 (
            .O(N__34200),
            .I(N__34197));
    LocalMux I__6634 (
            .O(N__34197),
            .I(N__34194));
    Odrv4 I__6633 (
            .O(N__34194),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    InMux I__6632 (
            .O(N__34191),
            .I(N__34188));
    LocalMux I__6631 (
            .O(N__34188),
            .I(N__34185));
    Odrv12 I__6630 (
            .O(N__34185),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__6629 (
            .O(N__34182),
            .I(N__34179));
    LocalMux I__6628 (
            .O(N__34179),
            .I(N__34176));
    Span4Mux_h I__6627 (
            .O(N__34176),
            .I(N__34173));
    Odrv4 I__6626 (
            .O(N__34173),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__6625 (
            .O(N__34170),
            .I(N__34167));
    LocalMux I__6624 (
            .O(N__34167),
            .I(N__34164));
    Span4Mux_h I__6623 (
            .O(N__34164),
            .I(N__34161));
    Odrv4 I__6622 (
            .O(N__34161),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__6621 (
            .O(N__34158),
            .I(N__34155));
    LocalMux I__6620 (
            .O(N__34155),
            .I(N__34152));
    Span4Mux_h I__6619 (
            .O(N__34152),
            .I(N__34149));
    Odrv4 I__6618 (
            .O(N__34149),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__6617 (
            .O(N__34146),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    CascadeMux I__6616 (
            .O(N__34143),
            .I(N__34139));
    InMux I__6615 (
            .O(N__34142),
            .I(N__34135));
    InMux I__6614 (
            .O(N__34139),
            .I(N__34130));
    InMux I__6613 (
            .O(N__34138),
            .I(N__34130));
    LocalMux I__6612 (
            .O(N__34135),
            .I(N__34127));
    LocalMux I__6611 (
            .O(N__34130),
            .I(N__34124));
    Span4Mux_v I__6610 (
            .O(N__34127),
            .I(N__34119));
    Span4Mux_h I__6609 (
            .O(N__34124),
            .I(N__34119));
    Odrv4 I__6608 (
            .O(N__34119),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__6607 (
            .O(N__34116),
            .I(N__34113));
    InMux I__6606 (
            .O(N__34113),
            .I(N__34110));
    LocalMux I__6605 (
            .O(N__34110),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    InMux I__6604 (
            .O(N__34107),
            .I(N__34104));
    LocalMux I__6603 (
            .O(N__34104),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    CascadeMux I__6602 (
            .O(N__34101),
            .I(elapsed_time_ns_1_RNII43T9_0_6_cascade_));
    CascadeMux I__6601 (
            .O(N__34098),
            .I(N__34095));
    InMux I__6600 (
            .O(N__34095),
            .I(N__34092));
    LocalMux I__6599 (
            .O(N__34092),
            .I(N__34089));
    Odrv4 I__6598 (
            .O(N__34089),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__6597 (
            .O(N__34086),
            .I(N__34082));
    InMux I__6596 (
            .O(N__34085),
            .I(N__34077));
    InMux I__6595 (
            .O(N__34082),
            .I(N__34077));
    LocalMux I__6594 (
            .O(N__34077),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    InMux I__6593 (
            .O(N__34074),
            .I(N__34071));
    LocalMux I__6592 (
            .O(N__34071),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__6591 (
            .O(N__34068),
            .I(N__34065));
    InMux I__6590 (
            .O(N__34065),
            .I(N__34062));
    LocalMux I__6589 (
            .O(N__34062),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__6588 (
            .O(N__34059),
            .I(N__34056));
    InMux I__6587 (
            .O(N__34056),
            .I(N__34053));
    LocalMux I__6586 (
            .O(N__34053),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__6585 (
            .O(N__34050),
            .I(N__34047));
    InMux I__6584 (
            .O(N__34047),
            .I(N__34044));
    LocalMux I__6583 (
            .O(N__34044),
            .I(N__34041));
    Odrv4 I__6582 (
            .O(N__34041),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__6581 (
            .O(N__34038),
            .I(N__34035));
    LocalMux I__6580 (
            .O(N__34035),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__6579 (
            .O(N__34032),
            .I(N__34029));
    InMux I__6578 (
            .O(N__34029),
            .I(N__34026));
    LocalMux I__6577 (
            .O(N__34026),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__6576 (
            .O(N__34023),
            .I(N__34020));
    LocalMux I__6575 (
            .O(N__34020),
            .I(N__34017));
    Span4Mux_v I__6574 (
            .O(N__34017),
            .I(N__34014));
    Odrv4 I__6573 (
            .O(N__34014),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__6572 (
            .O(N__34011),
            .I(N__34008));
    InMux I__6571 (
            .O(N__34008),
            .I(N__34005));
    LocalMux I__6570 (
            .O(N__34005),
            .I(N__34002));
    Odrv4 I__6569 (
            .O(N__34002),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__6568 (
            .O(N__33999),
            .I(N__33996));
    InMux I__6567 (
            .O(N__33996),
            .I(N__33993));
    LocalMux I__6566 (
            .O(N__33993),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__6565 (
            .O(N__33990),
            .I(N__33987));
    LocalMux I__6564 (
            .O(N__33987),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__6563 (
            .O(N__33984),
            .I(N__33981));
    InMux I__6562 (
            .O(N__33981),
            .I(N__33978));
    LocalMux I__6561 (
            .O(N__33978),
            .I(N__33975));
    Odrv4 I__6560 (
            .O(N__33975),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__6559 (
            .O(N__33972),
            .I(N__33969));
    InMux I__6558 (
            .O(N__33969),
            .I(N__33966));
    LocalMux I__6557 (
            .O(N__33966),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__6556 (
            .O(N__33963),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__6555 (
            .O(N__33960),
            .I(N__33954));
    InMux I__6554 (
            .O(N__33959),
            .I(N__33954));
    LocalMux I__6553 (
            .O(N__33954),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    CascadeMux I__6552 (
            .O(N__33951),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ));
    InMux I__6551 (
            .O(N__33948),
            .I(N__33945));
    LocalMux I__6550 (
            .O(N__33945),
            .I(N__33939));
    InMux I__6549 (
            .O(N__33944),
            .I(N__33932));
    InMux I__6548 (
            .O(N__33943),
            .I(N__33932));
    InMux I__6547 (
            .O(N__33942),
            .I(N__33932));
    Odrv4 I__6546 (
            .O(N__33939),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__6545 (
            .O(N__33932),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__6544 (
            .O(N__33927),
            .I(N__33924));
    InMux I__6543 (
            .O(N__33924),
            .I(N__33918));
    InMux I__6542 (
            .O(N__33923),
            .I(N__33918));
    LocalMux I__6541 (
            .O(N__33918),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__6540 (
            .O(N__33915),
            .I(N__33912));
    InMux I__6539 (
            .O(N__33912),
            .I(N__33909));
    LocalMux I__6538 (
            .O(N__33909),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__6537 (
            .O(N__33906),
            .I(N__33903));
    InMux I__6536 (
            .O(N__33903),
            .I(N__33900));
    LocalMux I__6535 (
            .O(N__33900),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__6534 (
            .O(N__33897),
            .I(N__33894));
    InMux I__6533 (
            .O(N__33894),
            .I(N__33891));
    LocalMux I__6532 (
            .O(N__33891),
            .I(N__33888));
    Odrv4 I__6531 (
            .O(N__33888),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__6530 (
            .O(N__33885),
            .I(N__33882));
    InMux I__6529 (
            .O(N__33882),
            .I(N__33879));
    LocalMux I__6528 (
            .O(N__33879),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__6527 (
            .O(N__33876),
            .I(N__33872));
    CascadeMux I__6526 (
            .O(N__33875),
            .I(N__33869));
    InMux I__6525 (
            .O(N__33872),
            .I(N__33861));
    InMux I__6524 (
            .O(N__33869),
            .I(N__33861));
    InMux I__6523 (
            .O(N__33868),
            .I(N__33861));
    LocalMux I__6522 (
            .O(N__33861),
            .I(\phase_controller_inst1.start_flagZ0 ));
    CascadeMux I__6521 (
            .O(N__33858),
            .I(N__33853));
    InMux I__6520 (
            .O(N__33857),
            .I(N__33850));
    InMux I__6519 (
            .O(N__33856),
            .I(N__33845));
    InMux I__6518 (
            .O(N__33853),
            .I(N__33845));
    LocalMux I__6517 (
            .O(N__33850),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6516 (
            .O(N__33845),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__6515 (
            .O(N__33840),
            .I(N__33837));
    LocalMux I__6514 (
            .O(N__33837),
            .I(\phase_controller_inst1.N_54_0 ));
    InMux I__6513 (
            .O(N__33834),
            .I(N__33830));
    InMux I__6512 (
            .O(N__33833),
            .I(N__33825));
    LocalMux I__6511 (
            .O(N__33830),
            .I(N__33822));
    InMux I__6510 (
            .O(N__33829),
            .I(N__33817));
    InMux I__6509 (
            .O(N__33828),
            .I(N__33817));
    LocalMux I__6508 (
            .O(N__33825),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__6507 (
            .O(N__33822),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__6506 (
            .O(N__33817),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__6505 (
            .O(N__33810),
            .I(N__33806));
    InMux I__6504 (
            .O(N__33809),
            .I(N__33803));
    LocalMux I__6503 (
            .O(N__33806),
            .I(N__33799));
    LocalMux I__6502 (
            .O(N__33803),
            .I(N__33796));
    InMux I__6501 (
            .O(N__33802),
            .I(N__33793));
    Span4Mux_h I__6500 (
            .O(N__33799),
            .I(N__33790));
    Span4Mux_h I__6499 (
            .O(N__33796),
            .I(N__33787));
    LocalMux I__6498 (
            .O(N__33793),
            .I(N__33784));
    Span4Mux_h I__6497 (
            .O(N__33790),
            .I(N__33781));
    Span4Mux_h I__6496 (
            .O(N__33787),
            .I(N__33778));
    IoSpan4Mux I__6495 (
            .O(N__33784),
            .I(N__33775));
    Odrv4 I__6494 (
            .O(N__33781),
            .I(il_max_comp1_c));
    Odrv4 I__6493 (
            .O(N__33778),
            .I(il_max_comp1_c));
    Odrv4 I__6492 (
            .O(N__33775),
            .I(il_max_comp1_c));
    CascadeMux I__6491 (
            .O(N__33768),
            .I(N__33765));
    InMux I__6490 (
            .O(N__33765),
            .I(N__33762));
    LocalMux I__6489 (
            .O(N__33762),
            .I(\phase_controller_inst2.state_ns_0_0_1 ));
    InMux I__6488 (
            .O(N__33759),
            .I(N__33756));
    LocalMux I__6487 (
            .O(N__33756),
            .I(N__33753));
    Sp12to4 I__6486 (
            .O(N__33753),
            .I(N__33750));
    Span12Mux_v I__6485 (
            .O(N__33750),
            .I(N__33744));
    InMux I__6484 (
            .O(N__33749),
            .I(N__33739));
    InMux I__6483 (
            .O(N__33748),
            .I(N__33739));
    InMux I__6482 (
            .O(N__33747),
            .I(N__33736));
    Odrv12 I__6481 (
            .O(N__33744),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__6480 (
            .O(N__33739),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__6479 (
            .O(N__33736),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    CascadeMux I__6478 (
            .O(N__33729),
            .I(N__33726));
    InMux I__6477 (
            .O(N__33726),
            .I(N__33721));
    InMux I__6476 (
            .O(N__33725),
            .I(N__33718));
    InMux I__6475 (
            .O(N__33724),
            .I(N__33715));
    LocalMux I__6474 (
            .O(N__33721),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__6473 (
            .O(N__33718),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__6472 (
            .O(N__33715),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__6471 (
            .O(N__33708),
            .I(N__33702));
    InMux I__6470 (
            .O(N__33707),
            .I(N__33702));
    LocalMux I__6469 (
            .O(N__33702),
            .I(\phase_controller_inst2.N_61 ));
    InMux I__6468 (
            .O(N__33699),
            .I(N__33659));
    InMux I__6467 (
            .O(N__33698),
            .I(N__33659));
    InMux I__6466 (
            .O(N__33697),
            .I(N__33659));
    InMux I__6465 (
            .O(N__33696),
            .I(N__33659));
    InMux I__6464 (
            .O(N__33695),
            .I(N__33650));
    InMux I__6463 (
            .O(N__33694),
            .I(N__33650));
    InMux I__6462 (
            .O(N__33693),
            .I(N__33650));
    InMux I__6461 (
            .O(N__33692),
            .I(N__33650));
    InMux I__6460 (
            .O(N__33691),
            .I(N__33643));
    InMux I__6459 (
            .O(N__33690),
            .I(N__33643));
    InMux I__6458 (
            .O(N__33689),
            .I(N__33643));
    InMux I__6457 (
            .O(N__33688),
            .I(N__33634));
    InMux I__6456 (
            .O(N__33687),
            .I(N__33634));
    InMux I__6455 (
            .O(N__33686),
            .I(N__33634));
    InMux I__6454 (
            .O(N__33685),
            .I(N__33634));
    IoInMux I__6453 (
            .O(N__33684),
            .I(N__33631));
    InMux I__6452 (
            .O(N__33683),
            .I(N__33628));
    InMux I__6451 (
            .O(N__33682),
            .I(N__33619));
    InMux I__6450 (
            .O(N__33681),
            .I(N__33619));
    InMux I__6449 (
            .O(N__33680),
            .I(N__33619));
    InMux I__6448 (
            .O(N__33679),
            .I(N__33619));
    InMux I__6447 (
            .O(N__33678),
            .I(N__33612));
    InMux I__6446 (
            .O(N__33677),
            .I(N__33612));
    InMux I__6445 (
            .O(N__33676),
            .I(N__33612));
    InMux I__6444 (
            .O(N__33675),
            .I(N__33603));
    InMux I__6443 (
            .O(N__33674),
            .I(N__33603));
    InMux I__6442 (
            .O(N__33673),
            .I(N__33603));
    InMux I__6441 (
            .O(N__33672),
            .I(N__33603));
    InMux I__6440 (
            .O(N__33671),
            .I(N__33594));
    InMux I__6439 (
            .O(N__33670),
            .I(N__33594));
    InMux I__6438 (
            .O(N__33669),
            .I(N__33594));
    InMux I__6437 (
            .O(N__33668),
            .I(N__33594));
    LocalMux I__6436 (
            .O(N__33659),
            .I(N__33589));
    LocalMux I__6435 (
            .O(N__33650),
            .I(N__33589));
    LocalMux I__6434 (
            .O(N__33643),
            .I(N__33586));
    LocalMux I__6433 (
            .O(N__33634),
            .I(N__33583));
    LocalMux I__6432 (
            .O(N__33631),
            .I(N__33580));
    LocalMux I__6431 (
            .O(N__33628),
            .I(N__33573));
    LocalMux I__6430 (
            .O(N__33619),
            .I(N__33573));
    LocalMux I__6429 (
            .O(N__33612),
            .I(N__33573));
    LocalMux I__6428 (
            .O(N__33603),
            .I(N__33562));
    LocalMux I__6427 (
            .O(N__33594),
            .I(N__33562));
    Span4Mux_h I__6426 (
            .O(N__33589),
            .I(N__33562));
    Span4Mux_v I__6425 (
            .O(N__33586),
            .I(N__33562));
    Span4Mux_v I__6424 (
            .O(N__33583),
            .I(N__33562));
    Span4Mux_s1_v I__6423 (
            .O(N__33580),
            .I(N__33559));
    Span4Mux_v I__6422 (
            .O(N__33573),
            .I(N__33552));
    Span4Mux_v I__6421 (
            .O(N__33562),
            .I(N__33552));
    Span4Mux_v I__6420 (
            .O(N__33559),
            .I(N__33552));
    Odrv4 I__6419 (
            .O(N__33552),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__6418 (
            .O(N__33549),
            .I(N__33546));
    LocalMux I__6417 (
            .O(N__33546),
            .I(\current_shift_inst.control_input_axb_27 ));
    ClkMux I__6416 (
            .O(N__33543),
            .I(N__33540));
    GlobalMux I__6415 (
            .O(N__33540),
            .I(N__33537));
    gio2CtrlBuf I__6414 (
            .O(N__33537),
            .I(delay_hc_input_c_g));
    IoInMux I__6413 (
            .O(N__33534),
            .I(N__33531));
    LocalMux I__6412 (
            .O(N__33531),
            .I(N__33528));
    IoSpan4Mux I__6411 (
            .O(N__33528),
            .I(N__33525));
    Span4Mux_s3_v I__6410 (
            .O(N__33525),
            .I(N__33522));
    Sp12to4 I__6409 (
            .O(N__33522),
            .I(N__33519));
    Odrv12 I__6408 (
            .O(N__33519),
            .I(s3_phy_c));
    IoInMux I__6407 (
            .O(N__33516),
            .I(N__33513));
    LocalMux I__6406 (
            .O(N__33513),
            .I(N__33510));
    Span4Mux_s0_v I__6405 (
            .O(N__33510),
            .I(N__33507));
    Odrv4 I__6404 (
            .O(N__33507),
            .I(GB_BUFFER_red_c_g_THRU_CO));
    InMux I__6403 (
            .O(N__33504),
            .I(N__33501));
    LocalMux I__6402 (
            .O(N__33501),
            .I(\phase_controller_inst1.state_ns_0_0_1 ));
    CascadeMux I__6401 (
            .O(N__33498),
            .I(N__33492));
    InMux I__6400 (
            .O(N__33497),
            .I(N__33489));
    InMux I__6399 (
            .O(N__33496),
            .I(N__33484));
    InMux I__6398 (
            .O(N__33495),
            .I(N__33484));
    InMux I__6397 (
            .O(N__33492),
            .I(N__33481));
    LocalMux I__6396 (
            .O(N__33489),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__6395 (
            .O(N__33484),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__6394 (
            .O(N__33481),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__6393 (
            .O(N__33474),
            .I(N__33470));
    InMux I__6392 (
            .O(N__33473),
            .I(N__33466));
    InMux I__6391 (
            .O(N__33470),
            .I(N__33463));
    InMux I__6390 (
            .O(N__33469),
            .I(N__33460));
    LocalMux I__6389 (
            .O(N__33466),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__6388 (
            .O(N__33463),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__6387 (
            .O(N__33460),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__6386 (
            .O(N__33453),
            .I(N__33444));
    InMux I__6385 (
            .O(N__33452),
            .I(N__33444));
    InMux I__6384 (
            .O(N__33451),
            .I(N__33444));
    LocalMux I__6383 (
            .O(N__33444),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    InMux I__6382 (
            .O(N__33441),
            .I(N__33438));
    LocalMux I__6381 (
            .O(N__33438),
            .I(\current_shift_inst.control_input_axb_14 ));
    InMux I__6380 (
            .O(N__33435),
            .I(N__33432));
    LocalMux I__6379 (
            .O(N__33432),
            .I(\current_shift_inst.control_input_axb_16 ));
    InMux I__6378 (
            .O(N__33429),
            .I(N__33426));
    LocalMux I__6377 (
            .O(N__33426),
            .I(\current_shift_inst.control_input_axb_18 ));
    InMux I__6376 (
            .O(N__33423),
            .I(N__33420));
    LocalMux I__6375 (
            .O(N__33420),
            .I(\current_shift_inst.control_input_axb_19 ));
    InMux I__6374 (
            .O(N__33417),
            .I(N__33414));
    LocalMux I__6373 (
            .O(N__33414),
            .I(\current_shift_inst.control_input_axb_20 ));
    InMux I__6372 (
            .O(N__33411),
            .I(N__33408));
    LocalMux I__6371 (
            .O(N__33408),
            .I(N__33405));
    Odrv4 I__6370 (
            .O(N__33405),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__6369 (
            .O(N__33402),
            .I(N__33399));
    LocalMux I__6368 (
            .O(N__33399),
            .I(\current_shift_inst.control_input_axb_23 ));
    InMux I__6367 (
            .O(N__33396),
            .I(N__33393));
    LocalMux I__6366 (
            .O(N__33393),
            .I(\current_shift_inst.control_input_axb_24 ));
    InMux I__6365 (
            .O(N__33390),
            .I(N__33387));
    LocalMux I__6364 (
            .O(N__33387),
            .I(\current_shift_inst.control_input_axb_25 ));
    InMux I__6363 (
            .O(N__33384),
            .I(N__33381));
    LocalMux I__6362 (
            .O(N__33381),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__6361 (
            .O(N__33378),
            .I(N__33375));
    LocalMux I__6360 (
            .O(N__33375),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__6359 (
            .O(N__33372),
            .I(N__33369));
    LocalMux I__6358 (
            .O(N__33369),
            .I(\current_shift_inst.control_input_axb_13 ));
    InMux I__6357 (
            .O(N__33366),
            .I(N__33363));
    LocalMux I__6356 (
            .O(N__33363),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__6355 (
            .O(N__33360),
            .I(N__33357));
    LocalMux I__6354 (
            .O(N__33357),
            .I(\current_shift_inst.control_input_axb_15 ));
    InMux I__6353 (
            .O(N__33354),
            .I(N__33350));
    InMux I__6352 (
            .O(N__33353),
            .I(N__33347));
    LocalMux I__6351 (
            .O(N__33350),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    LocalMux I__6350 (
            .O(N__33347),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CEMux I__6349 (
            .O(N__33342),
            .I(N__33306));
    CEMux I__6348 (
            .O(N__33341),
            .I(N__33306));
    CEMux I__6347 (
            .O(N__33340),
            .I(N__33306));
    CEMux I__6346 (
            .O(N__33339),
            .I(N__33306));
    CEMux I__6345 (
            .O(N__33338),
            .I(N__33306));
    CEMux I__6344 (
            .O(N__33337),
            .I(N__33306));
    CEMux I__6343 (
            .O(N__33336),
            .I(N__33306));
    CEMux I__6342 (
            .O(N__33335),
            .I(N__33306));
    CEMux I__6341 (
            .O(N__33334),
            .I(N__33306));
    CEMux I__6340 (
            .O(N__33333),
            .I(N__33306));
    CEMux I__6339 (
            .O(N__33332),
            .I(N__33306));
    CEMux I__6338 (
            .O(N__33331),
            .I(N__33306));
    GlobalMux I__6337 (
            .O(N__33306),
            .I(N__33303));
    gio2CtrlBuf I__6336 (
            .O(N__33303),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    InMux I__6335 (
            .O(N__33300),
            .I(N__33297));
    LocalMux I__6334 (
            .O(N__33297),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__6333 (
            .O(N__33294),
            .I(N__33290));
    InMux I__6332 (
            .O(N__33293),
            .I(N__33287));
    LocalMux I__6331 (
            .O(N__33290),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    LocalMux I__6330 (
            .O(N__33287),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    InMux I__6329 (
            .O(N__33282),
            .I(N__33277));
    InMux I__6328 (
            .O(N__33281),
            .I(N__33274));
    InMux I__6327 (
            .O(N__33280),
            .I(N__33271));
    LocalMux I__6326 (
            .O(N__33277),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__6325 (
            .O(N__33274),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__6324 (
            .O(N__33271),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    CascadeMux I__6323 (
            .O(N__33264),
            .I(N__33260));
    CascadeMux I__6322 (
            .O(N__33263),
            .I(N__33257));
    InMux I__6321 (
            .O(N__33260),
            .I(N__33254));
    InMux I__6320 (
            .O(N__33257),
            .I(N__33251));
    LocalMux I__6319 (
            .O(N__33254),
            .I(N__33246));
    LocalMux I__6318 (
            .O(N__33251),
            .I(N__33246));
    Span4Mux_v I__6317 (
            .O(N__33246),
            .I(N__33243));
    Odrv4 I__6316 (
            .O(N__33243),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    InMux I__6315 (
            .O(N__33240),
            .I(N__33235));
    InMux I__6314 (
            .O(N__33239),
            .I(N__33232));
    InMux I__6313 (
            .O(N__33238),
            .I(N__33229));
    LocalMux I__6312 (
            .O(N__33235),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__6311 (
            .O(N__33232),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__6310 (
            .O(N__33229),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__6309 (
            .O(N__33222),
            .I(N__33219));
    LocalMux I__6308 (
            .O(N__33219),
            .I(N__33216));
    Span4Mux_h I__6307 (
            .O(N__33216),
            .I(N__33213));
    Odrv4 I__6306 (
            .O(N__33213),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    InMux I__6305 (
            .O(N__33210),
            .I(N__33207));
    LocalMux I__6304 (
            .O(N__33207),
            .I(\current_shift_inst.control_input_axb_6 ));
    CascadeMux I__6303 (
            .O(N__33204),
            .I(N__33198));
    InMux I__6302 (
            .O(N__33203),
            .I(N__33195));
    InMux I__6301 (
            .O(N__33202),
            .I(N__33192));
    InMux I__6300 (
            .O(N__33201),
            .I(N__33189));
    InMux I__6299 (
            .O(N__33198),
            .I(N__33186));
    LocalMux I__6298 (
            .O(N__33195),
            .I(N__33183));
    LocalMux I__6297 (
            .O(N__33192),
            .I(N__33180));
    LocalMux I__6296 (
            .O(N__33189),
            .I(N__33175));
    LocalMux I__6295 (
            .O(N__33186),
            .I(N__33175));
    Span4Mux_v I__6294 (
            .O(N__33183),
            .I(N__33172));
    Span4Mux_v I__6293 (
            .O(N__33180),
            .I(N__33169));
    Span4Mux_v I__6292 (
            .O(N__33175),
            .I(N__33166));
    Odrv4 I__6291 (
            .O(N__33172),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__6290 (
            .O(N__33169),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__6289 (
            .O(N__33166),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__6288 (
            .O(N__33159),
            .I(N__33156));
    LocalMux I__6287 (
            .O(N__33156),
            .I(N__33152));
    InMux I__6286 (
            .O(N__33155),
            .I(N__33149));
    Span4Mux_v I__6285 (
            .O(N__33152),
            .I(N__33143));
    LocalMux I__6284 (
            .O(N__33149),
            .I(N__33143));
    InMux I__6283 (
            .O(N__33148),
            .I(N__33140));
    Span4Mux_h I__6282 (
            .O(N__33143),
            .I(N__33137));
    LocalMux I__6281 (
            .O(N__33140),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    Odrv4 I__6280 (
            .O(N__33137),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    CascadeMux I__6279 (
            .O(N__33132),
            .I(N__33129));
    InMux I__6278 (
            .O(N__33129),
            .I(N__33126));
    LocalMux I__6277 (
            .O(N__33126),
            .I(N__33123));
    Odrv4 I__6276 (
            .O(N__33123),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ));
    InMux I__6275 (
            .O(N__33120),
            .I(N__33114));
    InMux I__6274 (
            .O(N__33119),
            .I(N__33114));
    LocalMux I__6273 (
            .O(N__33114),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    CascadeMux I__6272 (
            .O(N__33111),
            .I(N__33108));
    InMux I__6271 (
            .O(N__33108),
            .I(N__33102));
    InMux I__6270 (
            .O(N__33107),
            .I(N__33102));
    LocalMux I__6269 (
            .O(N__33102),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    InMux I__6268 (
            .O(N__33099),
            .I(N__33096));
    LocalMux I__6267 (
            .O(N__33096),
            .I(N__33093));
    Span4Mux_h I__6266 (
            .O(N__33093),
            .I(N__33090));
    Odrv4 I__6265 (
            .O(N__33090),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    CascadeMux I__6264 (
            .O(N__33087),
            .I(N__33084));
    InMux I__6263 (
            .O(N__33084),
            .I(N__33081));
    LocalMux I__6262 (
            .O(N__33081),
            .I(N__33078));
    Span4Mux_v I__6261 (
            .O(N__33078),
            .I(N__33075));
    Odrv4 I__6260 (
            .O(N__33075),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    InMux I__6259 (
            .O(N__33072),
            .I(N__33069));
    LocalMux I__6258 (
            .O(N__33069),
            .I(N__33064));
    InMux I__6257 (
            .O(N__33068),
            .I(N__33061));
    InMux I__6256 (
            .O(N__33067),
            .I(N__33058));
    Span4Mux_h I__6255 (
            .O(N__33064),
            .I(N__33054));
    LocalMux I__6254 (
            .O(N__33061),
            .I(N__33051));
    LocalMux I__6253 (
            .O(N__33058),
            .I(N__33048));
    InMux I__6252 (
            .O(N__33057),
            .I(N__33045));
    Span4Mux_v I__6251 (
            .O(N__33054),
            .I(N__33042));
    Span4Mux_h I__6250 (
            .O(N__33051),
            .I(N__33037));
    Span4Mux_v I__6249 (
            .O(N__33048),
            .I(N__33037));
    LocalMux I__6248 (
            .O(N__33045),
            .I(N__33034));
    Odrv4 I__6247 (
            .O(N__33042),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__6246 (
            .O(N__33037),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv12 I__6245 (
            .O(N__33034),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__6244 (
            .O(N__33027),
            .I(N__33023));
    InMux I__6243 (
            .O(N__33026),
            .I(N__33019));
    LocalMux I__6242 (
            .O(N__33023),
            .I(N__33016));
    InMux I__6241 (
            .O(N__33022),
            .I(N__33013));
    LocalMux I__6240 (
            .O(N__33019),
            .I(N__33008));
    Span4Mux_v I__6239 (
            .O(N__33016),
            .I(N__33008));
    LocalMux I__6238 (
            .O(N__33013),
            .I(N__33005));
    Odrv4 I__6237 (
            .O(N__33008),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv4 I__6236 (
            .O(N__33005),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__6235 (
            .O(N__33000),
            .I(N__32995));
    InMux I__6234 (
            .O(N__32999),
            .I(N__32992));
    InMux I__6233 (
            .O(N__32998),
            .I(N__32989));
    LocalMux I__6232 (
            .O(N__32995),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__6231 (
            .O(N__32992),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__6230 (
            .O(N__32989),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__6229 (
            .O(N__32982),
            .I(N__32978));
    InMux I__6228 (
            .O(N__32981),
            .I(N__32975));
    LocalMux I__6227 (
            .O(N__32978),
            .I(N__32970));
    LocalMux I__6226 (
            .O(N__32975),
            .I(N__32970));
    Odrv12 I__6225 (
            .O(N__32970),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__6224 (
            .O(N__32967),
            .I(N__32963));
    CascadeMux I__6223 (
            .O(N__32966),
            .I(N__32959));
    InMux I__6222 (
            .O(N__32963),
            .I(N__32956));
    InMux I__6221 (
            .O(N__32962),
            .I(N__32953));
    InMux I__6220 (
            .O(N__32959),
            .I(N__32950));
    LocalMux I__6219 (
            .O(N__32956),
            .I(N__32947));
    LocalMux I__6218 (
            .O(N__32953),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__6217 (
            .O(N__32950),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__6216 (
            .O(N__32947),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__6215 (
            .O(N__32940),
            .I(N__32937));
    InMux I__6214 (
            .O(N__32937),
            .I(N__32934));
    LocalMux I__6213 (
            .O(N__32934),
            .I(N__32931));
    Span4Mux_h I__6212 (
            .O(N__32931),
            .I(N__32928));
    Span4Mux_h I__6211 (
            .O(N__32928),
            .I(N__32925));
    Odrv4 I__6210 (
            .O(N__32925),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    InMux I__6209 (
            .O(N__32922),
            .I(N__32919));
    LocalMux I__6208 (
            .O(N__32919),
            .I(N__32916));
    Span4Mux_v I__6207 (
            .O(N__32916),
            .I(N__32911));
    InMux I__6206 (
            .O(N__32915),
            .I(N__32906));
    InMux I__6205 (
            .O(N__32914),
            .I(N__32906));
    Sp12to4 I__6204 (
            .O(N__32911),
            .I(N__32901));
    LocalMux I__6203 (
            .O(N__32906),
            .I(N__32901));
    Span12Mux_h I__6202 (
            .O(N__32901),
            .I(N__32898));
    Odrv12 I__6201 (
            .O(N__32898),
            .I(il_max_comp2_c));
    InMux I__6200 (
            .O(N__32895),
            .I(N__32892));
    LocalMux I__6199 (
            .O(N__32892),
            .I(N__32889));
    Span4Mux_v I__6198 (
            .O(N__32889),
            .I(N__32884));
    InMux I__6197 (
            .O(N__32888),
            .I(N__32881));
    InMux I__6196 (
            .O(N__32887),
            .I(N__32878));
    Sp12to4 I__6195 (
            .O(N__32884),
            .I(N__32871));
    LocalMux I__6194 (
            .O(N__32881),
            .I(N__32871));
    LocalMux I__6193 (
            .O(N__32878),
            .I(N__32871));
    Span12Mux_h I__6192 (
            .O(N__32871),
            .I(N__32868));
    Odrv12 I__6191 (
            .O(N__32868),
            .I(il_min_comp2_c));
    InMux I__6190 (
            .O(N__32865),
            .I(N__32862));
    LocalMux I__6189 (
            .O(N__32862),
            .I(N__32859));
    Span4Mux_v I__6188 (
            .O(N__32859),
            .I(N__32855));
    InMux I__6187 (
            .O(N__32858),
            .I(N__32851));
    Sp12to4 I__6186 (
            .O(N__32855),
            .I(N__32848));
    InMux I__6185 (
            .O(N__32854),
            .I(N__32844));
    LocalMux I__6184 (
            .O(N__32851),
            .I(N__32839));
    Span12Mux_v I__6183 (
            .O(N__32848),
            .I(N__32839));
    InMux I__6182 (
            .O(N__32847),
            .I(N__32836));
    LocalMux I__6181 (
            .O(N__32844),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv12 I__6180 (
            .O(N__32839),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__6179 (
            .O(N__32836),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__6178 (
            .O(N__32829),
            .I(N__32824));
    InMux I__6177 (
            .O(N__32828),
            .I(N__32821));
    InMux I__6176 (
            .O(N__32827),
            .I(N__32818));
    LocalMux I__6175 (
            .O(N__32824),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__6174 (
            .O(N__32821),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__6173 (
            .O(N__32818),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__6172 (
            .O(N__32811),
            .I(N__32808));
    LocalMux I__6171 (
            .O(N__32808),
            .I(N__32805));
    Odrv4 I__6170 (
            .O(N__32805),
            .I(\phase_controller_inst2.N_54_0 ));
    CascadeMux I__6169 (
            .O(N__32802),
            .I(N__32798));
    CascadeMux I__6168 (
            .O(N__32801),
            .I(N__32793));
    InMux I__6167 (
            .O(N__32798),
            .I(N__32790));
    InMux I__6166 (
            .O(N__32797),
            .I(N__32785));
    InMux I__6165 (
            .O(N__32796),
            .I(N__32785));
    InMux I__6164 (
            .O(N__32793),
            .I(N__32782));
    LocalMux I__6163 (
            .O(N__32790),
            .I(N__32779));
    LocalMux I__6162 (
            .O(N__32785),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__6161 (
            .O(N__32782),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv4 I__6160 (
            .O(N__32779),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__6159 (
            .O(N__32772),
            .I(N__32767));
    CascadeMux I__6158 (
            .O(N__32771),
            .I(N__32764));
    InMux I__6157 (
            .O(N__32770),
            .I(N__32761));
    InMux I__6156 (
            .O(N__32767),
            .I(N__32758));
    InMux I__6155 (
            .O(N__32764),
            .I(N__32755));
    LocalMux I__6154 (
            .O(N__32761),
            .I(N__32752));
    LocalMux I__6153 (
            .O(N__32758),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__6152 (
            .O(N__32755),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__6151 (
            .O(N__32752),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__6150 (
            .O(N__32745),
            .I(N__32741));
    CascadeMux I__6149 (
            .O(N__32744),
            .I(N__32738));
    InMux I__6148 (
            .O(N__32741),
            .I(N__32734));
    InMux I__6147 (
            .O(N__32738),
            .I(N__32729));
    InMux I__6146 (
            .O(N__32737),
            .I(N__32729));
    LocalMux I__6145 (
            .O(N__32734),
            .I(N__32726));
    LocalMux I__6144 (
            .O(N__32729),
            .I(N__32723));
    Span4Mux_h I__6143 (
            .O(N__32726),
            .I(N__32720));
    Span4Mux_h I__6142 (
            .O(N__32723),
            .I(N__32717));
    Odrv4 I__6141 (
            .O(N__32720),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__6140 (
            .O(N__32717),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    CascadeMux I__6139 (
            .O(N__32712),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__6138 (
            .O(N__32709),
            .I(N__32706));
    LocalMux I__6137 (
            .O(N__32706),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__6136 (
            .O(N__32703),
            .I(N__32699));
    InMux I__6135 (
            .O(N__32702),
            .I(N__32696));
    LocalMux I__6134 (
            .O(N__32699),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__6133 (
            .O(N__32696),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    InMux I__6132 (
            .O(N__32691),
            .I(N__32688));
    LocalMux I__6131 (
            .O(N__32688),
            .I(N__32685));
    Span4Mux_v I__6130 (
            .O(N__32685),
            .I(N__32680));
    InMux I__6129 (
            .O(N__32684),
            .I(N__32677));
    InMux I__6128 (
            .O(N__32683),
            .I(N__32674));
    Span4Mux_h I__6127 (
            .O(N__32680),
            .I(N__32669));
    LocalMux I__6126 (
            .O(N__32677),
            .I(N__32669));
    LocalMux I__6125 (
            .O(N__32674),
            .I(N__32666));
    Sp12to4 I__6124 (
            .O(N__32669),
            .I(N__32663));
    Span4Mux_h I__6123 (
            .O(N__32666),
            .I(N__32659));
    Span12Mux_s10_v I__6122 (
            .O(N__32663),
            .I(N__32656));
    InMux I__6121 (
            .O(N__32662),
            .I(N__32653));
    Odrv4 I__6120 (
            .O(N__32659),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv12 I__6119 (
            .O(N__32656),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__6118 (
            .O(N__32653),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__6117 (
            .O(N__32646),
            .I(N__32643));
    LocalMux I__6116 (
            .O(N__32643),
            .I(N__32640));
    Span4Mux_h I__6115 (
            .O(N__32640),
            .I(N__32635));
    InMux I__6114 (
            .O(N__32639),
            .I(N__32632));
    InMux I__6113 (
            .O(N__32638),
            .I(N__32629));
    Span4Mux_v I__6112 (
            .O(N__32635),
            .I(N__32626));
    LocalMux I__6111 (
            .O(N__32632),
            .I(N__32623));
    LocalMux I__6110 (
            .O(N__32629),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__6109 (
            .O(N__32626),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv12 I__6108 (
            .O(N__32623),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__6107 (
            .O(N__32616),
            .I(N__32612));
    CascadeMux I__6106 (
            .O(N__32615),
            .I(N__32609));
    LocalMux I__6105 (
            .O(N__32612),
            .I(N__32606));
    InMux I__6104 (
            .O(N__32609),
            .I(N__32600));
    Span4Mux_s2_v I__6103 (
            .O(N__32606),
            .I(N__32597));
    InMux I__6102 (
            .O(N__32605),
            .I(N__32590));
    InMux I__6101 (
            .O(N__32604),
            .I(N__32590));
    InMux I__6100 (
            .O(N__32603),
            .I(N__32590));
    LocalMux I__6099 (
            .O(N__32600),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv4 I__6098 (
            .O(N__32597),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__6097 (
            .O(N__32590),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    CascadeMux I__6096 (
            .O(N__32583),
            .I(N__32579));
    InMux I__6095 (
            .O(N__32582),
            .I(N__32576));
    InMux I__6094 (
            .O(N__32579),
            .I(N__32572));
    LocalMux I__6093 (
            .O(N__32576),
            .I(N__32569));
    InMux I__6092 (
            .O(N__32575),
            .I(N__32566));
    LocalMux I__6091 (
            .O(N__32572),
            .I(N__32559));
    Span4Mux_h I__6090 (
            .O(N__32569),
            .I(N__32559));
    LocalMux I__6089 (
            .O(N__32566),
            .I(N__32559));
    Odrv4 I__6088 (
            .O(N__32559),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    CascadeMux I__6087 (
            .O(N__32556),
            .I(N__32552));
    InMux I__6086 (
            .O(N__32555),
            .I(N__32545));
    InMux I__6085 (
            .O(N__32552),
            .I(N__32545));
    InMux I__6084 (
            .O(N__32551),
            .I(N__32540));
    InMux I__6083 (
            .O(N__32550),
            .I(N__32540));
    LocalMux I__6082 (
            .O(N__32545),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__6081 (
            .O(N__32540),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__6080 (
            .O(N__32535),
            .I(N__32528));
    InMux I__6079 (
            .O(N__32534),
            .I(N__32528));
    InMux I__6078 (
            .O(N__32533),
            .I(N__32523));
    LocalMux I__6077 (
            .O(N__32528),
            .I(N__32520));
    InMux I__6076 (
            .O(N__32527),
            .I(N__32515));
    InMux I__6075 (
            .O(N__32526),
            .I(N__32515));
    LocalMux I__6074 (
            .O(N__32523),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__6073 (
            .O(N__32520),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__6072 (
            .O(N__32515),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__6071 (
            .O(N__32508),
            .I(N__32503));
    InMux I__6070 (
            .O(N__32507),
            .I(N__32500));
    InMux I__6069 (
            .O(N__32506),
            .I(N__32497));
    LocalMux I__6068 (
            .O(N__32503),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    LocalMux I__6067 (
            .O(N__32500),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    LocalMux I__6066 (
            .O(N__32497),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__6065 (
            .O(N__32490),
            .I(N__32487));
    LocalMux I__6064 (
            .O(N__32487),
            .I(N__32482));
    InMux I__6063 (
            .O(N__32486),
            .I(N__32479));
    InMux I__6062 (
            .O(N__32485),
            .I(N__32476));
    Span4Mux_h I__6061 (
            .O(N__32482),
            .I(N__32471));
    LocalMux I__6060 (
            .O(N__32479),
            .I(N__32471));
    LocalMux I__6059 (
            .O(N__32476),
            .I(N__32467));
    Span4Mux_h I__6058 (
            .O(N__32471),
            .I(N__32464));
    InMux I__6057 (
            .O(N__32470),
            .I(N__32461));
    Span12Mux_s11_v I__6056 (
            .O(N__32467),
            .I(N__32458));
    Span4Mux_v I__6055 (
            .O(N__32464),
            .I(N__32453));
    LocalMux I__6054 (
            .O(N__32461),
            .I(N__32453));
    Odrv12 I__6053 (
            .O(N__32458),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv4 I__6052 (
            .O(N__32453),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__6051 (
            .O(N__32448),
            .I(N__32445));
    LocalMux I__6050 (
            .O(N__32445),
            .I(N__32442));
    Odrv4 I__6049 (
            .O(N__32442),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ));
    InMux I__6048 (
            .O(N__32439),
            .I(\current_shift_inst.control_input_cry_25 ));
    InMux I__6047 (
            .O(N__32436),
            .I(N__32433));
    LocalMux I__6046 (
            .O(N__32433),
            .I(N__32430));
    Odrv4 I__6045 (
            .O(N__32430),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ));
    InMux I__6044 (
            .O(N__32427),
            .I(\current_shift_inst.control_input_cry_26 ));
    CascadeMux I__6043 (
            .O(N__32424),
            .I(N__32421));
    InMux I__6042 (
            .O(N__32421),
            .I(N__32418));
    LocalMux I__6041 (
            .O(N__32418),
            .I(N__32415));
    Odrv4 I__6040 (
            .O(N__32415),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ));
    InMux I__6039 (
            .O(N__32412),
            .I(\current_shift_inst.control_input_cry_27 ));
    CascadeMux I__6038 (
            .O(N__32409),
            .I(N__32406));
    InMux I__6037 (
            .O(N__32406),
            .I(N__32403));
    LocalMux I__6036 (
            .O(N__32403),
            .I(N__32400));
    Odrv4 I__6035 (
            .O(N__32400),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ));
    InMux I__6034 (
            .O(N__32397),
            .I(\current_shift_inst.control_input_cry_28 ));
    InMux I__6033 (
            .O(N__32394),
            .I(\current_shift_inst.control_input_cry_29 ));
    InMux I__6032 (
            .O(N__32391),
            .I(N__32388));
    LocalMux I__6031 (
            .O(N__32388),
            .I(N__32384));
    InMux I__6030 (
            .O(N__32387),
            .I(N__32381));
    Odrv4 I__6029 (
            .O(N__32384),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__6028 (
            .O(N__32381),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__6027 (
            .O(N__32376),
            .I(N__32373));
    LocalMux I__6026 (
            .O(N__32373),
            .I(\current_shift_inst.control_input_axb_26 ));
    InMux I__6025 (
            .O(N__32370),
            .I(N__32367));
    LocalMux I__6024 (
            .O(N__32367),
            .I(\current_shift_inst.control_input_axb_29 ));
    InMux I__6023 (
            .O(N__32364),
            .I(N__32361));
    LocalMux I__6022 (
            .O(N__32361),
            .I(N__32358));
    Odrv4 I__6021 (
            .O(N__32358),
            .I(\current_shift_inst.control_input_axb_17 ));
    IoInMux I__6020 (
            .O(N__32355),
            .I(N__32352));
    LocalMux I__6019 (
            .O(N__32352),
            .I(N__32349));
    IoSpan4Mux I__6018 (
            .O(N__32349),
            .I(N__32346));
    Span4Mux_s2_v I__6017 (
            .O(N__32346),
            .I(N__32343));
    Odrv4 I__6016 (
            .O(N__32343),
            .I(s4_phy_c));
    InMux I__6015 (
            .O(N__32340),
            .I(N__32337));
    LocalMux I__6014 (
            .O(N__32337),
            .I(N__32334));
    Odrv4 I__6013 (
            .O(N__32334),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    InMux I__6012 (
            .O(N__32331),
            .I(\current_shift_inst.control_input_cry_17 ));
    InMux I__6011 (
            .O(N__32328),
            .I(N__32325));
    LocalMux I__6010 (
            .O(N__32325),
            .I(N__32322));
    Odrv4 I__6009 (
            .O(N__32322),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__6008 (
            .O(N__32319),
            .I(\current_shift_inst.control_input_cry_18 ));
    CascadeMux I__6007 (
            .O(N__32316),
            .I(N__32313));
    InMux I__6006 (
            .O(N__32313),
            .I(N__32310));
    LocalMux I__6005 (
            .O(N__32310),
            .I(N__32307));
    Odrv4 I__6004 (
            .O(N__32307),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__6003 (
            .O(N__32304),
            .I(\current_shift_inst.control_input_cry_19 ));
    InMux I__6002 (
            .O(N__32301),
            .I(N__32298));
    LocalMux I__6001 (
            .O(N__32298),
            .I(N__32295));
    Odrv4 I__6000 (
            .O(N__32295),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__5999 (
            .O(N__32292),
            .I(\current_shift_inst.control_input_cry_20 ));
    CascadeMux I__5998 (
            .O(N__32289),
            .I(N__32286));
    InMux I__5997 (
            .O(N__32286),
            .I(N__32283));
    LocalMux I__5996 (
            .O(N__32283),
            .I(N__32280));
    Odrv4 I__5995 (
            .O(N__32280),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__5994 (
            .O(N__32277),
            .I(\current_shift_inst.control_input_cry_21 ));
    CascadeMux I__5993 (
            .O(N__32274),
            .I(N__32271));
    InMux I__5992 (
            .O(N__32271),
            .I(N__32268));
    LocalMux I__5991 (
            .O(N__32268),
            .I(N__32265));
    Odrv4 I__5990 (
            .O(N__32265),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__5989 (
            .O(N__32262),
            .I(\current_shift_inst.control_input_cry_22 ));
    InMux I__5988 (
            .O(N__32259),
            .I(N__32256));
    LocalMux I__5987 (
            .O(N__32256),
            .I(N__32253));
    Odrv4 I__5986 (
            .O(N__32253),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__5985 (
            .O(N__32250),
            .I(bfn_11_16_0_));
    InMux I__5984 (
            .O(N__32247),
            .I(N__32244));
    LocalMux I__5983 (
            .O(N__32244),
            .I(N__32241));
    Odrv4 I__5982 (
            .O(N__32241),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__5981 (
            .O(N__32238),
            .I(\current_shift_inst.control_input_cry_24 ));
    CascadeMux I__5980 (
            .O(N__32235),
            .I(N__32232));
    InMux I__5979 (
            .O(N__32232),
            .I(N__32229));
    LocalMux I__5978 (
            .O(N__32229),
            .I(N__32226));
    Odrv4 I__5977 (
            .O(N__32226),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__5976 (
            .O(N__32223),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__5975 (
            .O(N__32220),
            .I(N__32217));
    LocalMux I__5974 (
            .O(N__32217),
            .I(N__32214));
    Odrv4 I__5973 (
            .O(N__32214),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__5972 (
            .O(N__32211),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__5971 (
            .O(N__32208),
            .I(N__32205));
    LocalMux I__5970 (
            .O(N__32205),
            .I(N__32202));
    Odrv4 I__5969 (
            .O(N__32202),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__5968 (
            .O(N__32199),
            .I(\current_shift_inst.control_input_cry_11 ));
    CascadeMux I__5967 (
            .O(N__32196),
            .I(N__32193));
    InMux I__5966 (
            .O(N__32193),
            .I(N__32190));
    LocalMux I__5965 (
            .O(N__32190),
            .I(N__32187));
    Odrv4 I__5964 (
            .O(N__32187),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__5963 (
            .O(N__32184),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__5962 (
            .O(N__32181),
            .I(N__32178));
    LocalMux I__5961 (
            .O(N__32178),
            .I(N__32175));
    Odrv4 I__5960 (
            .O(N__32175),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__5959 (
            .O(N__32172),
            .I(\current_shift_inst.control_input_cry_13 ));
    CascadeMux I__5958 (
            .O(N__32169),
            .I(N__32166));
    InMux I__5957 (
            .O(N__32166),
            .I(N__32163));
    LocalMux I__5956 (
            .O(N__32163),
            .I(N__32160));
    Odrv4 I__5955 (
            .O(N__32160),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__5954 (
            .O(N__32157),
            .I(\current_shift_inst.control_input_cry_14 ));
    InMux I__5953 (
            .O(N__32154),
            .I(N__32151));
    LocalMux I__5952 (
            .O(N__32151),
            .I(N__32148));
    Odrv4 I__5951 (
            .O(N__32148),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__5950 (
            .O(N__32145),
            .I(bfn_11_15_0_));
    CascadeMux I__5949 (
            .O(N__32142),
            .I(N__32139));
    InMux I__5948 (
            .O(N__32139),
            .I(N__32136));
    LocalMux I__5947 (
            .O(N__32136),
            .I(N__32133));
    Odrv4 I__5946 (
            .O(N__32133),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__5945 (
            .O(N__32130),
            .I(\current_shift_inst.control_input_cry_16 ));
    InMux I__5944 (
            .O(N__32127),
            .I(N__32124));
    LocalMux I__5943 (
            .O(N__32124),
            .I(N__32121));
    Odrv4 I__5942 (
            .O(N__32121),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__5941 (
            .O(N__32118),
            .I(\current_shift_inst.control_input_cry_0 ));
    CascadeMux I__5940 (
            .O(N__32115),
            .I(N__32112));
    InMux I__5939 (
            .O(N__32112),
            .I(N__32109));
    LocalMux I__5938 (
            .O(N__32109),
            .I(N__32106));
    Odrv4 I__5937 (
            .O(N__32106),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__5936 (
            .O(N__32103),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__5935 (
            .O(N__32100),
            .I(N__32097));
    LocalMux I__5934 (
            .O(N__32097),
            .I(N__32094));
    Odrv4 I__5933 (
            .O(N__32094),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__5932 (
            .O(N__32091),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__5931 (
            .O(N__32088),
            .I(N__32085));
    LocalMux I__5930 (
            .O(N__32085),
            .I(N__32082));
    Odrv4 I__5929 (
            .O(N__32082),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__5928 (
            .O(N__32079),
            .I(\current_shift_inst.control_input_cry_3 ));
    CascadeMux I__5927 (
            .O(N__32076),
            .I(N__32073));
    InMux I__5926 (
            .O(N__32073),
            .I(N__32070));
    LocalMux I__5925 (
            .O(N__32070),
            .I(N__32067));
    Odrv4 I__5924 (
            .O(N__32067),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__5923 (
            .O(N__32064),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__5922 (
            .O(N__32061),
            .I(N__32058));
    LocalMux I__5921 (
            .O(N__32058),
            .I(N__32055));
    Odrv4 I__5920 (
            .O(N__32055),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__5919 (
            .O(N__32052),
            .I(\current_shift_inst.control_input_cry_5 ));
    CascadeMux I__5918 (
            .O(N__32049),
            .I(N__32046));
    InMux I__5917 (
            .O(N__32046),
            .I(N__32043));
    LocalMux I__5916 (
            .O(N__32043),
            .I(N__32040));
    Odrv4 I__5915 (
            .O(N__32040),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__5914 (
            .O(N__32037),
            .I(\current_shift_inst.control_input_cry_6 ));
    CascadeMux I__5913 (
            .O(N__32034),
            .I(N__32031));
    InMux I__5912 (
            .O(N__32031),
            .I(N__32028));
    LocalMux I__5911 (
            .O(N__32028),
            .I(N__32025));
    Odrv4 I__5910 (
            .O(N__32025),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__5909 (
            .O(N__32022),
            .I(bfn_11_14_0_));
    InMux I__5908 (
            .O(N__32019),
            .I(N__32016));
    LocalMux I__5907 (
            .O(N__32016),
            .I(N__32013));
    Odrv4 I__5906 (
            .O(N__32013),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__5905 (
            .O(N__32010),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__5904 (
            .O(N__32007),
            .I(N__32002));
    InMux I__5903 (
            .O(N__32006),
            .I(N__31997));
    InMux I__5902 (
            .O(N__32005),
            .I(N__31997));
    LocalMux I__5901 (
            .O(N__32002),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__5900 (
            .O(N__31997),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__5899 (
            .O(N__31992),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    CascadeMux I__5898 (
            .O(N__31989),
            .I(N__31985));
    InMux I__5897 (
            .O(N__31988),
            .I(N__31979));
    InMux I__5896 (
            .O(N__31985),
            .I(N__31979));
    InMux I__5895 (
            .O(N__31984),
            .I(N__31976));
    LocalMux I__5894 (
            .O(N__31979),
            .I(N__31973));
    LocalMux I__5893 (
            .O(N__31976),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__5892 (
            .O(N__31973),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__5891 (
            .O(N__31968),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__5890 (
            .O(N__31965),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__5889 (
            .O(N__31962),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    CascadeMux I__5888 (
            .O(N__31959),
            .I(N__31954));
    InMux I__5887 (
            .O(N__31958),
            .I(N__31951));
    InMux I__5886 (
            .O(N__31957),
            .I(N__31946));
    InMux I__5885 (
            .O(N__31954),
            .I(N__31946));
    LocalMux I__5884 (
            .O(N__31951),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__5883 (
            .O(N__31946),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__5882 (
            .O(N__31941),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__5881 (
            .O(N__31938),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__5880 (
            .O(N__31935),
            .I(N__31930));
    InMux I__5879 (
            .O(N__31934),
            .I(N__31925));
    InMux I__5878 (
            .O(N__31933),
            .I(N__31925));
    LocalMux I__5877 (
            .O(N__31930),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__5876 (
            .O(N__31925),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    CascadeMux I__5875 (
            .O(N__31920),
            .I(N__31915));
    InMux I__5874 (
            .O(N__31919),
            .I(N__31912));
    InMux I__5873 (
            .O(N__31918),
            .I(N__31909));
    InMux I__5872 (
            .O(N__31915),
            .I(N__31906));
    LocalMux I__5871 (
            .O(N__31912),
            .I(\current_shift_inst.N_1263_i ));
    LocalMux I__5870 (
            .O(N__31909),
            .I(\current_shift_inst.N_1263_i ));
    LocalMux I__5869 (
            .O(N__31906),
            .I(\current_shift_inst.N_1263_i ));
    InMux I__5868 (
            .O(N__31899),
            .I(N__31896));
    LocalMux I__5867 (
            .O(N__31896),
            .I(N__31893));
    Odrv4 I__5866 (
            .O(N__31893),
            .I(\current_shift_inst.control_input_1 ));
    InMux I__5865 (
            .O(N__31890),
            .I(bfn_11_10_0_));
    CascadeMux I__5864 (
            .O(N__31887),
            .I(N__31883));
    InMux I__5863 (
            .O(N__31886),
            .I(N__31877));
    InMux I__5862 (
            .O(N__31883),
            .I(N__31877));
    InMux I__5861 (
            .O(N__31882),
            .I(N__31874));
    LocalMux I__5860 (
            .O(N__31877),
            .I(N__31871));
    LocalMux I__5859 (
            .O(N__31874),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__5858 (
            .O(N__31871),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__5857 (
            .O(N__31866),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__5856 (
            .O(N__31863),
            .I(N__31856));
    InMux I__5855 (
            .O(N__31862),
            .I(N__31856));
    InMux I__5854 (
            .O(N__31861),
            .I(N__31853));
    LocalMux I__5853 (
            .O(N__31856),
            .I(N__31850));
    LocalMux I__5852 (
            .O(N__31853),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__5851 (
            .O(N__31850),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__5850 (
            .O(N__31845),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__5849 (
            .O(N__31842),
            .I(N__31835));
    InMux I__5848 (
            .O(N__31841),
            .I(N__31835));
    InMux I__5847 (
            .O(N__31840),
            .I(N__31832));
    LocalMux I__5846 (
            .O(N__31835),
            .I(N__31829));
    LocalMux I__5845 (
            .O(N__31832),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__5844 (
            .O(N__31829),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__5843 (
            .O(N__31824),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    CascadeMux I__5842 (
            .O(N__31821),
            .I(N__31817));
    InMux I__5841 (
            .O(N__31820),
            .I(N__31811));
    InMux I__5840 (
            .O(N__31817),
            .I(N__31811));
    InMux I__5839 (
            .O(N__31816),
            .I(N__31808));
    LocalMux I__5838 (
            .O(N__31811),
            .I(N__31805));
    LocalMux I__5837 (
            .O(N__31808),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__5836 (
            .O(N__31805),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__5835 (
            .O(N__31800),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__5834 (
            .O(N__31797),
            .I(N__31793));
    InMux I__5833 (
            .O(N__31796),
            .I(N__31787));
    InMux I__5832 (
            .O(N__31793),
            .I(N__31787));
    InMux I__5831 (
            .O(N__31792),
            .I(N__31784));
    LocalMux I__5830 (
            .O(N__31787),
            .I(N__31781));
    LocalMux I__5829 (
            .O(N__31784),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv12 I__5828 (
            .O(N__31781),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__5827 (
            .O(N__31776),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__5826 (
            .O(N__31773),
            .I(N__31766));
    InMux I__5825 (
            .O(N__31772),
            .I(N__31766));
    InMux I__5824 (
            .O(N__31771),
            .I(N__31763));
    LocalMux I__5823 (
            .O(N__31766),
            .I(N__31760));
    LocalMux I__5822 (
            .O(N__31763),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv12 I__5821 (
            .O(N__31760),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__5820 (
            .O(N__31755),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__5819 (
            .O(N__31752),
            .I(N__31746));
    InMux I__5818 (
            .O(N__31751),
            .I(N__31746));
    LocalMux I__5817 (
            .O(N__31746),
            .I(N__31742));
    InMux I__5816 (
            .O(N__31745),
            .I(N__31739));
    Span4Mux_h I__5815 (
            .O(N__31742),
            .I(N__31736));
    LocalMux I__5814 (
            .O(N__31739),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__5813 (
            .O(N__31736),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__5812 (
            .O(N__31731),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    CascadeMux I__5811 (
            .O(N__31728),
            .I(N__31724));
    InMux I__5810 (
            .O(N__31727),
            .I(N__31719));
    InMux I__5809 (
            .O(N__31724),
            .I(N__31719));
    LocalMux I__5808 (
            .O(N__31719),
            .I(N__31715));
    InMux I__5807 (
            .O(N__31718),
            .I(N__31712));
    Span4Mux_h I__5806 (
            .O(N__31715),
            .I(N__31709));
    LocalMux I__5805 (
            .O(N__31712),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__5804 (
            .O(N__31709),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__5803 (
            .O(N__31704),
            .I(bfn_11_11_0_));
    InMux I__5802 (
            .O(N__31701),
            .I(N__31697));
    InMux I__5801 (
            .O(N__31700),
            .I(N__31694));
    LocalMux I__5800 (
            .O(N__31697),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__5799 (
            .O(N__31694),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__5798 (
            .O(N__31689),
            .I(bfn_11_9_0_));
    InMux I__5797 (
            .O(N__31686),
            .I(N__31682));
    InMux I__5796 (
            .O(N__31685),
            .I(N__31679));
    LocalMux I__5795 (
            .O(N__31682),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__5794 (
            .O(N__31679),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__5793 (
            .O(N__31674),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__5792 (
            .O(N__31671),
            .I(N__31667));
    InMux I__5791 (
            .O(N__31670),
            .I(N__31664));
    LocalMux I__5790 (
            .O(N__31667),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__5789 (
            .O(N__31664),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__5788 (
            .O(N__31659),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__5787 (
            .O(N__31656),
            .I(N__31652));
    InMux I__5786 (
            .O(N__31655),
            .I(N__31649));
    LocalMux I__5785 (
            .O(N__31652),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__5784 (
            .O(N__31649),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__5783 (
            .O(N__31644),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__5782 (
            .O(N__31641),
            .I(N__31637));
    InMux I__5781 (
            .O(N__31640),
            .I(N__31634));
    LocalMux I__5780 (
            .O(N__31637),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__5779 (
            .O(N__31634),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__5778 (
            .O(N__31629),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__5777 (
            .O(N__31626),
            .I(N__31622));
    InMux I__5776 (
            .O(N__31625),
            .I(N__31619));
    LocalMux I__5775 (
            .O(N__31622),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__5774 (
            .O(N__31619),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__5773 (
            .O(N__31614),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__5772 (
            .O(N__31611),
            .I(N__31607));
    InMux I__5771 (
            .O(N__31610),
            .I(N__31604));
    LocalMux I__5770 (
            .O(N__31607),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__5769 (
            .O(N__31604),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__5768 (
            .O(N__31599),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__5767 (
            .O(N__31596),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__5766 (
            .O(N__31593),
            .I(N__31588));
    InMux I__5765 (
            .O(N__31592),
            .I(N__31583));
    InMux I__5764 (
            .O(N__31591),
            .I(N__31583));
    LocalMux I__5763 (
            .O(N__31588),
            .I(N__31580));
    LocalMux I__5762 (
            .O(N__31583),
            .I(N__31577));
    Span4Mux_v I__5761 (
            .O(N__31580),
            .I(N__31571));
    Span4Mux_v I__5760 (
            .O(N__31577),
            .I(N__31571));
    InMux I__5759 (
            .O(N__31576),
            .I(N__31568));
    Span4Mux_h I__5758 (
            .O(N__31571),
            .I(N__31563));
    LocalMux I__5757 (
            .O(N__31568),
            .I(N__31563));
    Odrv4 I__5756 (
            .O(N__31563),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__5755 (
            .O(N__31560),
            .I(N__31556));
    InMux I__5754 (
            .O(N__31559),
            .I(N__31553));
    LocalMux I__5753 (
            .O(N__31556),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    LocalMux I__5752 (
            .O(N__31553),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    CascadeMux I__5751 (
            .O(N__31548),
            .I(N__31545));
    InMux I__5750 (
            .O(N__31545),
            .I(N__31542));
    LocalMux I__5749 (
            .O(N__31542),
            .I(N__31539));
    Odrv4 I__5748 (
            .O(N__31539),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    InMux I__5747 (
            .O(N__31536),
            .I(N__31532));
    InMux I__5746 (
            .O(N__31535),
            .I(N__31529));
    LocalMux I__5745 (
            .O(N__31532),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__5744 (
            .O(N__31529),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__5743 (
            .O(N__31524),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__5742 (
            .O(N__31521),
            .I(N__31517));
    InMux I__5741 (
            .O(N__31520),
            .I(N__31514));
    LocalMux I__5740 (
            .O(N__31517),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__5739 (
            .O(N__31514),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__5738 (
            .O(N__31509),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__5737 (
            .O(N__31506),
            .I(N__31502));
    InMux I__5736 (
            .O(N__31505),
            .I(N__31499));
    LocalMux I__5735 (
            .O(N__31502),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__5734 (
            .O(N__31499),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__5733 (
            .O(N__31494),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__5732 (
            .O(N__31491),
            .I(N__31487));
    InMux I__5731 (
            .O(N__31490),
            .I(N__31484));
    LocalMux I__5730 (
            .O(N__31487),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__5729 (
            .O(N__31484),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__5728 (
            .O(N__31479),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__5727 (
            .O(N__31476),
            .I(N__31472));
    InMux I__5726 (
            .O(N__31475),
            .I(N__31469));
    LocalMux I__5725 (
            .O(N__31472),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__5724 (
            .O(N__31469),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__5723 (
            .O(N__31464),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__5722 (
            .O(N__31461),
            .I(N__31457));
    InMux I__5721 (
            .O(N__31460),
            .I(N__31454));
    LocalMux I__5720 (
            .O(N__31457),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__5719 (
            .O(N__31454),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__5718 (
            .O(N__31449),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__5717 (
            .O(N__31446),
            .I(N__31442));
    InMux I__5716 (
            .O(N__31445),
            .I(N__31439));
    LocalMux I__5715 (
            .O(N__31442),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__5714 (
            .O(N__31439),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__5713 (
            .O(N__31434),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__5712 (
            .O(N__31431),
            .I(N__31427));
    InMux I__5711 (
            .O(N__31430),
            .I(N__31424));
    LocalMux I__5710 (
            .O(N__31427),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    LocalMux I__5709 (
            .O(N__31424),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__5708 (
            .O(N__31419),
            .I(N__31415));
    InMux I__5707 (
            .O(N__31418),
            .I(N__31411));
    LocalMux I__5706 (
            .O(N__31415),
            .I(N__31408));
    InMux I__5705 (
            .O(N__31414),
            .I(N__31405));
    LocalMux I__5704 (
            .O(N__31411),
            .I(N__31402));
    Span4Mux_s2_v I__5703 (
            .O(N__31408),
            .I(N__31397));
    LocalMux I__5702 (
            .O(N__31405),
            .I(N__31397));
    Span4Mux_h I__5701 (
            .O(N__31402),
            .I(N__31392));
    Span4Mux_v I__5700 (
            .O(N__31397),
            .I(N__31392));
    Span4Mux_v I__5699 (
            .O(N__31392),
            .I(N__31388));
    InMux I__5698 (
            .O(N__31391),
            .I(N__31385));
    Odrv4 I__5697 (
            .O(N__31388),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__5696 (
            .O(N__31385),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__5695 (
            .O(N__31380),
            .I(N__31377));
    LocalMux I__5694 (
            .O(N__31377),
            .I(N__31372));
    InMux I__5693 (
            .O(N__31376),
            .I(N__31369));
    InMux I__5692 (
            .O(N__31375),
            .I(N__31366));
    Span4Mux_v I__5691 (
            .O(N__31372),
            .I(N__31361));
    LocalMux I__5690 (
            .O(N__31369),
            .I(N__31361));
    LocalMux I__5689 (
            .O(N__31366),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv4 I__5688 (
            .O(N__31361),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__5687 (
            .O(N__31356),
            .I(N__31352));
    InMux I__5686 (
            .O(N__31355),
            .I(N__31349));
    LocalMux I__5685 (
            .O(N__31352),
            .I(N__31345));
    LocalMux I__5684 (
            .O(N__31349),
            .I(N__31342));
    InMux I__5683 (
            .O(N__31348),
            .I(N__31339));
    Span4Mux_h I__5682 (
            .O(N__31345),
            .I(N__31333));
    Span4Mux_h I__5681 (
            .O(N__31342),
            .I(N__31333));
    LocalMux I__5680 (
            .O(N__31339),
            .I(N__31330));
    InMux I__5679 (
            .O(N__31338),
            .I(N__31327));
    Span4Mux_v I__5678 (
            .O(N__31333),
            .I(N__31324));
    Span4Mux_v I__5677 (
            .O(N__31330),
            .I(N__31321));
    LocalMux I__5676 (
            .O(N__31327),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv4 I__5675 (
            .O(N__31324),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv4 I__5674 (
            .O(N__31321),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__5673 (
            .O(N__31314),
            .I(N__31311));
    LocalMux I__5672 (
            .O(N__31311),
            .I(N__31308));
    Span4Mux_h I__5671 (
            .O(N__31308),
            .I(N__31303));
    InMux I__5670 (
            .O(N__31307),
            .I(N__31300));
    InMux I__5669 (
            .O(N__31306),
            .I(N__31297));
    Span4Mux_v I__5668 (
            .O(N__31303),
            .I(N__31294));
    LocalMux I__5667 (
            .O(N__31300),
            .I(N__31291));
    LocalMux I__5666 (
            .O(N__31297),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    Odrv4 I__5665 (
            .O(N__31294),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    Odrv12 I__5664 (
            .O(N__31291),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    CascadeMux I__5663 (
            .O(N__31284),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_));
    InMux I__5662 (
            .O(N__31281),
            .I(N__31278));
    LocalMux I__5661 (
            .O(N__31278),
            .I(N__31275));
    Span4Mux_s1_v I__5660 (
            .O(N__31275),
            .I(N__31272));
    Span4Mux_v I__5659 (
            .O(N__31272),
            .I(N__31269));
    Odrv4 I__5658 (
            .O(N__31269),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    CEMux I__5657 (
            .O(N__31266),
            .I(N__31260));
    CEMux I__5656 (
            .O(N__31265),
            .I(N__31257));
    CEMux I__5655 (
            .O(N__31264),
            .I(N__31251));
    CEMux I__5654 (
            .O(N__31263),
            .I(N__31245));
    LocalMux I__5653 (
            .O(N__31260),
            .I(N__31240));
    LocalMux I__5652 (
            .O(N__31257),
            .I(N__31240));
    CEMux I__5651 (
            .O(N__31256),
            .I(N__31220));
    CEMux I__5650 (
            .O(N__31255),
            .I(N__31208));
    CEMux I__5649 (
            .O(N__31254),
            .I(N__31205));
    LocalMux I__5648 (
            .O(N__31251),
            .I(N__31202));
    CEMux I__5647 (
            .O(N__31250),
            .I(N__31196));
    CEMux I__5646 (
            .O(N__31249),
            .I(N__31193));
    CEMux I__5645 (
            .O(N__31248),
            .I(N__31190));
    LocalMux I__5644 (
            .O(N__31245),
            .I(N__31185));
    Span4Mux_h I__5643 (
            .O(N__31240),
            .I(N__31185));
    InMux I__5642 (
            .O(N__31239),
            .I(N__31178));
    InMux I__5641 (
            .O(N__31238),
            .I(N__31178));
    InMux I__5640 (
            .O(N__31237),
            .I(N__31178));
    InMux I__5639 (
            .O(N__31236),
            .I(N__31169));
    InMux I__5638 (
            .O(N__31235),
            .I(N__31169));
    InMux I__5637 (
            .O(N__31234),
            .I(N__31169));
    InMux I__5636 (
            .O(N__31233),
            .I(N__31169));
    InMux I__5635 (
            .O(N__31232),
            .I(N__31166));
    InMux I__5634 (
            .O(N__31231),
            .I(N__31157));
    InMux I__5633 (
            .O(N__31230),
            .I(N__31157));
    InMux I__5632 (
            .O(N__31229),
            .I(N__31157));
    InMux I__5631 (
            .O(N__31228),
            .I(N__31157));
    InMux I__5630 (
            .O(N__31227),
            .I(N__31148));
    InMux I__5629 (
            .O(N__31226),
            .I(N__31148));
    InMux I__5628 (
            .O(N__31225),
            .I(N__31148));
    InMux I__5627 (
            .O(N__31224),
            .I(N__31148));
    CEMux I__5626 (
            .O(N__31223),
            .I(N__31145));
    LocalMux I__5625 (
            .O(N__31220),
            .I(N__31142));
    InMux I__5624 (
            .O(N__31219),
            .I(N__31133));
    InMux I__5623 (
            .O(N__31218),
            .I(N__31133));
    InMux I__5622 (
            .O(N__31217),
            .I(N__31133));
    InMux I__5621 (
            .O(N__31216),
            .I(N__31133));
    InMux I__5620 (
            .O(N__31215),
            .I(N__31124));
    InMux I__5619 (
            .O(N__31214),
            .I(N__31124));
    InMux I__5618 (
            .O(N__31213),
            .I(N__31124));
    InMux I__5617 (
            .O(N__31212),
            .I(N__31124));
    CEMux I__5616 (
            .O(N__31211),
            .I(N__31114));
    LocalMux I__5615 (
            .O(N__31208),
            .I(N__31109));
    LocalMux I__5614 (
            .O(N__31205),
            .I(N__31109));
    Span4Mux_h I__5613 (
            .O(N__31202),
            .I(N__31106));
    CEMux I__5612 (
            .O(N__31201),
            .I(N__31103));
    CEMux I__5611 (
            .O(N__31200),
            .I(N__31100));
    CEMux I__5610 (
            .O(N__31199),
            .I(N__31097));
    LocalMux I__5609 (
            .O(N__31196),
            .I(N__31092));
    LocalMux I__5608 (
            .O(N__31193),
            .I(N__31092));
    LocalMux I__5607 (
            .O(N__31190),
            .I(N__31083));
    Span4Mux_v I__5606 (
            .O(N__31185),
            .I(N__31083));
    LocalMux I__5605 (
            .O(N__31178),
            .I(N__31083));
    LocalMux I__5604 (
            .O(N__31169),
            .I(N__31083));
    LocalMux I__5603 (
            .O(N__31166),
            .I(N__31080));
    LocalMux I__5602 (
            .O(N__31157),
            .I(N__31075));
    LocalMux I__5601 (
            .O(N__31148),
            .I(N__31075));
    LocalMux I__5600 (
            .O(N__31145),
            .I(N__31068));
    Span4Mux_s3_v I__5599 (
            .O(N__31142),
            .I(N__31068));
    LocalMux I__5598 (
            .O(N__31133),
            .I(N__31068));
    LocalMux I__5597 (
            .O(N__31124),
            .I(N__31065));
    InMux I__5596 (
            .O(N__31123),
            .I(N__31058));
    InMux I__5595 (
            .O(N__31122),
            .I(N__31058));
    InMux I__5594 (
            .O(N__31121),
            .I(N__31058));
    InMux I__5593 (
            .O(N__31120),
            .I(N__31049));
    InMux I__5592 (
            .O(N__31119),
            .I(N__31049));
    InMux I__5591 (
            .O(N__31118),
            .I(N__31049));
    InMux I__5590 (
            .O(N__31117),
            .I(N__31049));
    LocalMux I__5589 (
            .O(N__31114),
            .I(N__31038));
    Span4Mux_v I__5588 (
            .O(N__31109),
            .I(N__31038));
    Span4Mux_h I__5587 (
            .O(N__31106),
            .I(N__31038));
    LocalMux I__5586 (
            .O(N__31103),
            .I(N__31038));
    LocalMux I__5585 (
            .O(N__31100),
            .I(N__31038));
    LocalMux I__5584 (
            .O(N__31097),
            .I(N__31031));
    Span4Mux_h I__5583 (
            .O(N__31092),
            .I(N__31031));
    Span4Mux_h I__5582 (
            .O(N__31083),
            .I(N__31031));
    Span4Mux_h I__5581 (
            .O(N__31080),
            .I(N__31026));
    Span4Mux_h I__5580 (
            .O(N__31075),
            .I(N__31026));
    Span4Mux_h I__5579 (
            .O(N__31068),
            .I(N__31021));
    Span4Mux_h I__5578 (
            .O(N__31065),
            .I(N__31021));
    LocalMux I__5577 (
            .O(N__31058),
            .I(N__31014));
    LocalMux I__5576 (
            .O(N__31049),
            .I(N__31014));
    Span4Mux_v I__5575 (
            .O(N__31038),
            .I(N__31014));
    Odrv4 I__5574 (
            .O(N__31031),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__5573 (
            .O(N__31026),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__5572 (
            .O(N__31021),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__5571 (
            .O(N__31014),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__5570 (
            .O(N__31005),
            .I(N__31001));
    InMux I__5569 (
            .O(N__31004),
            .I(N__30997));
    LocalMux I__5568 (
            .O(N__31001),
            .I(N__30994));
    InMux I__5567 (
            .O(N__31000),
            .I(N__30991));
    LocalMux I__5566 (
            .O(N__30997),
            .I(N__30988));
    Span4Mux_h I__5565 (
            .O(N__30994),
            .I(N__30985));
    LocalMux I__5564 (
            .O(N__30991),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv4 I__5563 (
            .O(N__30988),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv4 I__5562 (
            .O(N__30985),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__5561 (
            .O(N__30978),
            .I(N__30974));
    InMux I__5560 (
            .O(N__30977),
            .I(N__30971));
    LocalMux I__5559 (
            .O(N__30974),
            .I(N__30967));
    LocalMux I__5558 (
            .O(N__30971),
            .I(N__30964));
    InMux I__5557 (
            .O(N__30970),
            .I(N__30961));
    Span4Mux_h I__5556 (
            .O(N__30967),
            .I(N__30953));
    Span4Mux_v I__5555 (
            .O(N__30964),
            .I(N__30953));
    LocalMux I__5554 (
            .O(N__30961),
            .I(N__30953));
    InMux I__5553 (
            .O(N__30960),
            .I(N__30950));
    Odrv4 I__5552 (
            .O(N__30953),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__5551 (
            .O(N__30950),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__5550 (
            .O(N__30945),
            .I(N__30942));
    LocalMux I__5549 (
            .O(N__30942),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__5548 (
            .O(N__30939),
            .I(N__30935));
    InMux I__5547 (
            .O(N__30938),
            .I(N__30930));
    InMux I__5546 (
            .O(N__30935),
            .I(N__30930));
    LocalMux I__5545 (
            .O(N__30930),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    InMux I__5544 (
            .O(N__30927),
            .I(N__30924));
    LocalMux I__5543 (
            .O(N__30924),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    InMux I__5542 (
            .O(N__30921),
            .I(N__30917));
    InMux I__5541 (
            .O(N__30920),
            .I(N__30913));
    LocalMux I__5540 (
            .O(N__30917),
            .I(N__30910));
    InMux I__5539 (
            .O(N__30916),
            .I(N__30907));
    LocalMux I__5538 (
            .O(N__30913),
            .I(N__30904));
    Span4Mux_h I__5537 (
            .O(N__30910),
            .I(N__30901));
    LocalMux I__5536 (
            .O(N__30907),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    Odrv12 I__5535 (
            .O(N__30904),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    Odrv4 I__5534 (
            .O(N__30901),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    InMux I__5533 (
            .O(N__30894),
            .I(N__30890));
    InMux I__5532 (
            .O(N__30893),
            .I(N__30886));
    LocalMux I__5531 (
            .O(N__30890),
            .I(N__30882));
    InMux I__5530 (
            .O(N__30889),
            .I(N__30879));
    LocalMux I__5529 (
            .O(N__30886),
            .I(N__30876));
    InMux I__5528 (
            .O(N__30885),
            .I(N__30873));
    Span4Mux_h I__5527 (
            .O(N__30882),
            .I(N__30868));
    LocalMux I__5526 (
            .O(N__30879),
            .I(N__30868));
    Sp12to4 I__5525 (
            .O(N__30876),
            .I(N__30863));
    LocalMux I__5524 (
            .O(N__30873),
            .I(N__30863));
    Odrv4 I__5523 (
            .O(N__30868),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv12 I__5522 (
            .O(N__30863),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__5521 (
            .O(N__30858),
            .I(N__30852));
    InMux I__5520 (
            .O(N__30857),
            .I(N__30852));
    LocalMux I__5519 (
            .O(N__30852),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__5518 (
            .O(N__30849),
            .I(N__30846));
    InMux I__5517 (
            .O(N__30846),
            .I(N__30843));
    LocalMux I__5516 (
            .O(N__30843),
            .I(N__30840));
    Odrv12 I__5515 (
            .O(N__30840),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    InMux I__5514 (
            .O(N__30837),
            .I(N__30831));
    InMux I__5513 (
            .O(N__30836),
            .I(N__30831));
    LocalMux I__5512 (
            .O(N__30831),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__5511 (
            .O(N__30828),
            .I(N__30825));
    InMux I__5510 (
            .O(N__30825),
            .I(N__30819));
    InMux I__5509 (
            .O(N__30824),
            .I(N__30819));
    LocalMux I__5508 (
            .O(N__30819),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__5507 (
            .O(N__30816),
            .I(N__30813));
    LocalMux I__5506 (
            .O(N__30813),
            .I(N__30810));
    Odrv4 I__5505 (
            .O(N__30810),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    InMux I__5504 (
            .O(N__30807),
            .I(N__30804));
    LocalMux I__5503 (
            .O(N__30804),
            .I(N__30800));
    InMux I__5502 (
            .O(N__30803),
            .I(N__30797));
    Span4Mux_v I__5501 (
            .O(N__30800),
            .I(N__30794));
    LocalMux I__5500 (
            .O(N__30797),
            .I(N__30791));
    Sp12to4 I__5499 (
            .O(N__30794),
            .I(N__30788));
    Span12Mux_v I__5498 (
            .O(N__30791),
            .I(N__30785));
    Span12Mux_s10_h I__5497 (
            .O(N__30788),
            .I(N__30782));
    Odrv12 I__5496 (
            .O(N__30785),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv12 I__5495 (
            .O(N__30782),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__5494 (
            .O(N__30777),
            .I(N__30774));
    LocalMux I__5493 (
            .O(N__30774),
            .I(N__30770));
    InMux I__5492 (
            .O(N__30773),
            .I(N__30766));
    Span4Mux_v I__5491 (
            .O(N__30770),
            .I(N__30763));
    InMux I__5490 (
            .O(N__30769),
            .I(N__30760));
    LocalMux I__5489 (
            .O(N__30766),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__5488 (
            .O(N__30763),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    LocalMux I__5487 (
            .O(N__30760),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__5486 (
            .O(N__30753),
            .I(N__30748));
    InMux I__5485 (
            .O(N__30752),
            .I(N__30745));
    InMux I__5484 (
            .O(N__30751),
            .I(N__30741));
    LocalMux I__5483 (
            .O(N__30748),
            .I(N__30736));
    LocalMux I__5482 (
            .O(N__30745),
            .I(N__30736));
    InMux I__5481 (
            .O(N__30744),
            .I(N__30733));
    LocalMux I__5480 (
            .O(N__30741),
            .I(N__30730));
    Span4Mux_v I__5479 (
            .O(N__30736),
            .I(N__30727));
    LocalMux I__5478 (
            .O(N__30733),
            .I(N__30724));
    Odrv4 I__5477 (
            .O(N__30730),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__5476 (
            .O(N__30727),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv12 I__5475 (
            .O(N__30724),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__5474 (
            .O(N__30717),
            .I(N__30714));
    LocalMux I__5473 (
            .O(N__30714),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ));
    InMux I__5472 (
            .O(N__30711),
            .I(N__30708));
    LocalMux I__5471 (
            .O(N__30708),
            .I(N__30705));
    Span4Mux_v I__5470 (
            .O(N__30705),
            .I(N__30702));
    Sp12to4 I__5469 (
            .O(N__30702),
            .I(N__30699));
    Span12Mux_h I__5468 (
            .O(N__30699),
            .I(N__30696));
    Odrv12 I__5467 (
            .O(N__30696),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__5466 (
            .O(N__30693),
            .I(N__30690));
    LocalMux I__5465 (
            .O(N__30690),
            .I(N__30687));
    Span4Mux_h I__5464 (
            .O(N__30687),
            .I(N__30684));
    Span4Mux_h I__5463 (
            .O(N__30684),
            .I(N__30681));
    Odrv4 I__5462 (
            .O(N__30681),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__5461 (
            .O(N__30678),
            .I(N__30675));
    LocalMux I__5460 (
            .O(N__30675),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    CascadeMux I__5459 (
            .O(N__30672),
            .I(N__30669));
    InMux I__5458 (
            .O(N__30669),
            .I(N__30666));
    LocalMux I__5457 (
            .O(N__30666),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    InMux I__5456 (
            .O(N__30663),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__5455 (
            .O(N__30660),
            .I(N__30657));
    InMux I__5454 (
            .O(N__30657),
            .I(N__30654));
    LocalMux I__5453 (
            .O(N__30654),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    CascadeMux I__5452 (
            .O(N__30651),
            .I(N__30647));
    InMux I__5451 (
            .O(N__30650),
            .I(N__30642));
    InMux I__5450 (
            .O(N__30647),
            .I(N__30642));
    LocalMux I__5449 (
            .O(N__30642),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    InMux I__5448 (
            .O(N__30639),
            .I(N__30636));
    LocalMux I__5447 (
            .O(N__30636),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    InMux I__5446 (
            .O(N__30633),
            .I(N__30628));
    InMux I__5445 (
            .O(N__30632),
            .I(N__30625));
    InMux I__5444 (
            .O(N__30631),
            .I(N__30622));
    LocalMux I__5443 (
            .O(N__30628),
            .I(N__30619));
    LocalMux I__5442 (
            .O(N__30625),
            .I(N__30616));
    LocalMux I__5441 (
            .O(N__30622),
            .I(N__30611));
    Span4Mux_v I__5440 (
            .O(N__30619),
            .I(N__30611));
    Odrv12 I__5439 (
            .O(N__30616),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    Odrv4 I__5438 (
            .O(N__30611),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    InMux I__5437 (
            .O(N__30606),
            .I(N__30601));
    CascadeMux I__5436 (
            .O(N__30605),
            .I(N__30598));
    InMux I__5435 (
            .O(N__30604),
            .I(N__30594));
    LocalMux I__5434 (
            .O(N__30601),
            .I(N__30591));
    InMux I__5433 (
            .O(N__30598),
            .I(N__30588));
    InMux I__5432 (
            .O(N__30597),
            .I(N__30585));
    LocalMux I__5431 (
            .O(N__30594),
            .I(N__30582));
    Span4Mux_v I__5430 (
            .O(N__30591),
            .I(N__30579));
    LocalMux I__5429 (
            .O(N__30588),
            .I(N__30576));
    LocalMux I__5428 (
            .O(N__30585),
            .I(N__30573));
    Span4Mux_h I__5427 (
            .O(N__30582),
            .I(N__30566));
    Span4Mux_v I__5426 (
            .O(N__30579),
            .I(N__30566));
    Span4Mux_v I__5425 (
            .O(N__30576),
            .I(N__30566));
    Odrv12 I__5424 (
            .O(N__30573),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__5423 (
            .O(N__30566),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__5422 (
            .O(N__30561),
            .I(N__30555));
    InMux I__5421 (
            .O(N__30560),
            .I(N__30555));
    LocalMux I__5420 (
            .O(N__30555),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    CascadeMux I__5419 (
            .O(N__30552),
            .I(N__30549));
    InMux I__5418 (
            .O(N__30549),
            .I(N__30546));
    LocalMux I__5417 (
            .O(N__30546),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    CascadeMux I__5416 (
            .O(N__30543),
            .I(N__30540));
    InMux I__5415 (
            .O(N__30540),
            .I(N__30537));
    LocalMux I__5414 (
            .O(N__30537),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    InMux I__5413 (
            .O(N__30534),
            .I(N__30531));
    LocalMux I__5412 (
            .O(N__30531),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__5411 (
            .O(N__30528),
            .I(N__30525));
    LocalMux I__5410 (
            .O(N__30525),
            .I(N__30522));
    Odrv4 I__5409 (
            .O(N__30522),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__5408 (
            .O(N__30519),
            .I(N__30516));
    InMux I__5407 (
            .O(N__30516),
            .I(N__30513));
    LocalMux I__5406 (
            .O(N__30513),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__5405 (
            .O(N__30510),
            .I(N__30507));
    LocalMux I__5404 (
            .O(N__30507),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__5403 (
            .O(N__30504),
            .I(N__30501));
    LocalMux I__5402 (
            .O(N__30501),
            .I(N__30498));
    Span4Mux_h I__5401 (
            .O(N__30498),
            .I(N__30495));
    Span4Mux_h I__5400 (
            .O(N__30495),
            .I(N__30492));
    Odrv4 I__5399 (
            .O(N__30492),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__5398 (
            .O(N__30489),
            .I(N__30486));
    InMux I__5397 (
            .O(N__30486),
            .I(N__30483));
    LocalMux I__5396 (
            .O(N__30483),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__5395 (
            .O(N__30480),
            .I(N__30477));
    LocalMux I__5394 (
            .O(N__30477),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    CascadeMux I__5393 (
            .O(N__30474),
            .I(N__30471));
    InMux I__5392 (
            .O(N__30471),
            .I(N__30468));
    LocalMux I__5391 (
            .O(N__30468),
            .I(N__30465));
    Odrv4 I__5390 (
            .O(N__30465),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    InMux I__5389 (
            .O(N__30462),
            .I(N__30459));
    LocalMux I__5388 (
            .O(N__30459),
            .I(N__30456));
    Odrv4 I__5387 (
            .O(N__30456),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    CascadeMux I__5386 (
            .O(N__30453),
            .I(N__30450));
    InMux I__5385 (
            .O(N__30450),
            .I(N__30447));
    LocalMux I__5384 (
            .O(N__30447),
            .I(N__30444));
    Odrv4 I__5383 (
            .O(N__30444),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__5382 (
            .O(N__30441),
            .I(N__30438));
    LocalMux I__5381 (
            .O(N__30438),
            .I(N__30435));
    Odrv4 I__5380 (
            .O(N__30435),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__5379 (
            .O(N__30432),
            .I(N__30429));
    InMux I__5378 (
            .O(N__30429),
            .I(N__30426));
    LocalMux I__5377 (
            .O(N__30426),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__5376 (
            .O(N__30423),
            .I(N__30420));
    LocalMux I__5375 (
            .O(N__30420),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__5374 (
            .O(N__30417),
            .I(N__30414));
    InMux I__5373 (
            .O(N__30414),
            .I(N__30411));
    LocalMux I__5372 (
            .O(N__30411),
            .I(N__30408));
    Odrv4 I__5371 (
            .O(N__30408),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__5370 (
            .O(N__30405),
            .I(N__30402));
    LocalMux I__5369 (
            .O(N__30402),
            .I(N__30399));
    Odrv4 I__5368 (
            .O(N__30399),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__5367 (
            .O(N__30396),
            .I(N__30393));
    InMux I__5366 (
            .O(N__30393),
            .I(N__30390));
    LocalMux I__5365 (
            .O(N__30390),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__5364 (
            .O(N__30387),
            .I(N__30384));
    LocalMux I__5363 (
            .O(N__30384),
            .I(N__30381));
    Span4Mux_v I__5362 (
            .O(N__30381),
            .I(N__30378));
    Odrv4 I__5361 (
            .O(N__30378),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__5360 (
            .O(N__30375),
            .I(N__30372));
    InMux I__5359 (
            .O(N__30372),
            .I(N__30369));
    LocalMux I__5358 (
            .O(N__30369),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__5357 (
            .O(N__30366),
            .I(N__30363));
    InMux I__5356 (
            .O(N__30363),
            .I(N__30360));
    LocalMux I__5355 (
            .O(N__30360),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__5354 (
            .O(N__30357),
            .I(N__30354));
    LocalMux I__5353 (
            .O(N__30354),
            .I(N__30351));
    Odrv4 I__5352 (
            .O(N__30351),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__5351 (
            .O(N__30348),
            .I(N__30345));
    InMux I__5350 (
            .O(N__30345),
            .I(N__30342));
    LocalMux I__5349 (
            .O(N__30342),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__5348 (
            .O(N__30339),
            .I(N__30336));
    LocalMux I__5347 (
            .O(N__30336),
            .I(N__30333));
    Odrv4 I__5346 (
            .O(N__30333),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__5345 (
            .O(N__30330),
            .I(N__30327));
    InMux I__5344 (
            .O(N__30327),
            .I(N__30324));
    LocalMux I__5343 (
            .O(N__30324),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__5342 (
            .O(N__30321),
            .I(N__30318));
    LocalMux I__5341 (
            .O(N__30318),
            .I(N__30315));
    Odrv4 I__5340 (
            .O(N__30315),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__5339 (
            .O(N__30312),
            .I(N__30309));
    InMux I__5338 (
            .O(N__30309),
            .I(N__30306));
    LocalMux I__5337 (
            .O(N__30306),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__5336 (
            .O(N__30303),
            .I(N__30300));
    LocalMux I__5335 (
            .O(N__30300),
            .I(N__30295));
    InMux I__5334 (
            .O(N__30299),
            .I(N__30292));
    InMux I__5333 (
            .O(N__30298),
            .I(N__30289));
    Span4Mux_s3_v I__5332 (
            .O(N__30295),
            .I(N__30284));
    LocalMux I__5331 (
            .O(N__30292),
            .I(N__30284));
    LocalMux I__5330 (
            .O(N__30289),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    Odrv4 I__5329 (
            .O(N__30284),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__5328 (
            .O(N__30279),
            .I(N__30275));
    InMux I__5327 (
            .O(N__30278),
            .I(N__30272));
    LocalMux I__5326 (
            .O(N__30275),
            .I(N__30268));
    LocalMux I__5325 (
            .O(N__30272),
            .I(N__30265));
    InMux I__5324 (
            .O(N__30271),
            .I(N__30261));
    Span4Mux_v I__5323 (
            .O(N__30268),
            .I(N__30256));
    Span4Mux_v I__5322 (
            .O(N__30265),
            .I(N__30256));
    CascadeMux I__5321 (
            .O(N__30264),
            .I(N__30253));
    LocalMux I__5320 (
            .O(N__30261),
            .I(N__30250));
    Span4Mux_v I__5319 (
            .O(N__30256),
            .I(N__30247));
    InMux I__5318 (
            .O(N__30253),
            .I(N__30244));
    Span12Mux_h I__5317 (
            .O(N__30250),
            .I(N__30241));
    Sp12to4 I__5316 (
            .O(N__30247),
            .I(N__30238));
    LocalMux I__5315 (
            .O(N__30244),
            .I(N__30235));
    Odrv12 I__5314 (
            .O(N__30241),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv12 I__5313 (
            .O(N__30238),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__5312 (
            .O(N__30235),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__5311 (
            .O(N__30228),
            .I(N__30224));
    InMux I__5310 (
            .O(N__30227),
            .I(N__30220));
    LocalMux I__5309 (
            .O(N__30224),
            .I(N__30217));
    InMux I__5308 (
            .O(N__30223),
            .I(N__30214));
    LocalMux I__5307 (
            .O(N__30220),
            .I(N__30210));
    Span4Mux_s2_v I__5306 (
            .O(N__30217),
            .I(N__30205));
    LocalMux I__5305 (
            .O(N__30214),
            .I(N__30205));
    InMux I__5304 (
            .O(N__30213),
            .I(N__30202));
    Span4Mux_h I__5303 (
            .O(N__30210),
            .I(N__30197));
    Span4Mux_v I__5302 (
            .O(N__30205),
            .I(N__30197));
    LocalMux I__5301 (
            .O(N__30202),
            .I(N__30194));
    Odrv4 I__5300 (
            .O(N__30197),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__5299 (
            .O(N__30194),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__5298 (
            .O(N__30189),
            .I(N__30186));
    LocalMux I__5297 (
            .O(N__30186),
            .I(N__30181));
    InMux I__5296 (
            .O(N__30185),
            .I(N__30178));
    InMux I__5295 (
            .O(N__30184),
            .I(N__30175));
    Span4Mux_h I__5294 (
            .O(N__30181),
            .I(N__30172));
    LocalMux I__5293 (
            .O(N__30178),
            .I(N__30169));
    LocalMux I__5292 (
            .O(N__30175),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv4 I__5291 (
            .O(N__30172),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv4 I__5290 (
            .O(N__30169),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__5289 (
            .O(N__30162),
            .I(N__30158));
    InMux I__5288 (
            .O(N__30161),
            .I(N__30155));
    LocalMux I__5287 (
            .O(N__30158),
            .I(N__30149));
    LocalMux I__5286 (
            .O(N__30155),
            .I(N__30149));
    InMux I__5285 (
            .O(N__30154),
            .I(N__30146));
    Sp12to4 I__5284 (
            .O(N__30149),
            .I(N__30140));
    LocalMux I__5283 (
            .O(N__30146),
            .I(N__30140));
    InMux I__5282 (
            .O(N__30145),
            .I(N__30137));
    Span12Mux_s10_v I__5281 (
            .O(N__30140),
            .I(N__30134));
    LocalMux I__5280 (
            .O(N__30137),
            .I(N__30131));
    Odrv12 I__5279 (
            .O(N__30134),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv12 I__5278 (
            .O(N__30131),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__5277 (
            .O(N__30126),
            .I(N__30122));
    InMux I__5276 (
            .O(N__30125),
            .I(N__30118));
    LocalMux I__5275 (
            .O(N__30122),
            .I(N__30115));
    InMux I__5274 (
            .O(N__30121),
            .I(N__30112));
    LocalMux I__5273 (
            .O(N__30118),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    Odrv4 I__5272 (
            .O(N__30115),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    LocalMux I__5271 (
            .O(N__30112),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    InMux I__5270 (
            .O(N__30105),
            .I(N__30100));
    InMux I__5269 (
            .O(N__30104),
            .I(N__30097));
    InMux I__5268 (
            .O(N__30103),
            .I(N__30094));
    LocalMux I__5267 (
            .O(N__30100),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__5266 (
            .O(N__30097),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__5265 (
            .O(N__30094),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__5264 (
            .O(N__30087),
            .I(N__30084));
    LocalMux I__5263 (
            .O(N__30084),
            .I(N__30080));
    InMux I__5262 (
            .O(N__30083),
            .I(N__30077));
    Span4Mux_h I__5261 (
            .O(N__30080),
            .I(N__30072));
    LocalMux I__5260 (
            .O(N__30077),
            .I(N__30069));
    InMux I__5259 (
            .O(N__30076),
            .I(N__30064));
    InMux I__5258 (
            .O(N__30075),
            .I(N__30064));
    Span4Mux_v I__5257 (
            .O(N__30072),
            .I(N__30061));
    Span4Mux_h I__5256 (
            .O(N__30069),
            .I(N__30058));
    LocalMux I__5255 (
            .O(N__30064),
            .I(N__30055));
    Odrv4 I__5254 (
            .O(N__30061),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    Odrv4 I__5253 (
            .O(N__30058),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    Odrv12 I__5252 (
            .O(N__30055),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    CascadeMux I__5251 (
            .O(N__30048),
            .I(N__30045));
    InMux I__5250 (
            .O(N__30045),
            .I(N__30042));
    LocalMux I__5249 (
            .O(N__30042),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    InMux I__5248 (
            .O(N__30039),
            .I(N__30036));
    LocalMux I__5247 (
            .O(N__30036),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__5246 (
            .O(N__30033),
            .I(N__30030));
    InMux I__5245 (
            .O(N__30030),
            .I(N__30027));
    LocalMux I__5244 (
            .O(N__30027),
            .I(N__30024));
    Odrv4 I__5243 (
            .O(N__30024),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    InMux I__5242 (
            .O(N__30021),
            .I(N__30018));
    LocalMux I__5241 (
            .O(N__30018),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__5240 (
            .O(N__30015),
            .I(N__30012));
    InMux I__5239 (
            .O(N__30012),
            .I(N__30009));
    LocalMux I__5238 (
            .O(N__30009),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    InMux I__5237 (
            .O(N__30006),
            .I(N__30003));
    LocalMux I__5236 (
            .O(N__30003),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__5235 (
            .O(N__30000),
            .I(N__29997));
    LocalMux I__5234 (
            .O(N__29997),
            .I(N__29993));
    InMux I__5233 (
            .O(N__29996),
            .I(N__29990));
    Odrv4 I__5232 (
            .O(N__29993),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__5231 (
            .O(N__29990),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__5230 (
            .O(N__29985),
            .I(N__29982));
    InMux I__5229 (
            .O(N__29982),
            .I(N__29979));
    LocalMux I__5228 (
            .O(N__29979),
            .I(N__29976));
    Odrv4 I__5227 (
            .O(N__29976),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ));
    InMux I__5226 (
            .O(N__29973),
            .I(N__29970));
    LocalMux I__5225 (
            .O(N__29970),
            .I(N__29967));
    Span12Mux_s10_h I__5224 (
            .O(N__29967),
            .I(N__29964));
    Odrv12 I__5223 (
            .O(N__29964),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__5222 (
            .O(N__29961),
            .I(N__29958));
    LocalMux I__5221 (
            .O(N__29958),
            .I(N__29955));
    Span4Mux_h I__5220 (
            .O(N__29955),
            .I(N__29952));
    Odrv4 I__5219 (
            .O(N__29952),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__5218 (
            .O(N__29949),
            .I(N__29943));
    InMux I__5217 (
            .O(N__29948),
            .I(N__29943));
    LocalMux I__5216 (
            .O(N__29943),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__5215 (
            .O(N__29940),
            .I(N__29935));
    InMux I__5214 (
            .O(N__29939),
            .I(N__29932));
    InMux I__5213 (
            .O(N__29938),
            .I(N__29927));
    InMux I__5212 (
            .O(N__29935),
            .I(N__29927));
    LocalMux I__5211 (
            .O(N__29932),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__5210 (
            .O(N__29927),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__5209 (
            .O(N__29922),
            .I(N__29918));
    InMux I__5208 (
            .O(N__29921),
            .I(N__29914));
    InMux I__5207 (
            .O(N__29918),
            .I(N__29911));
    InMux I__5206 (
            .O(N__29917),
            .I(N__29908));
    LocalMux I__5205 (
            .O(N__29914),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__5204 (
            .O(N__29911),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__5203 (
            .O(N__29908),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__5202 (
            .O(N__29901),
            .I(N__29898));
    InMux I__5201 (
            .O(N__29898),
            .I(N__29895));
    LocalMux I__5200 (
            .O(N__29895),
            .I(N__29892));
    Span4Mux_h I__5199 (
            .O(N__29892),
            .I(N__29889));
    Odrv4 I__5198 (
            .O(N__29889),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    InMux I__5197 (
            .O(N__29886),
            .I(N__29882));
    InMux I__5196 (
            .O(N__29885),
            .I(N__29879));
    LocalMux I__5195 (
            .O(N__29882),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    LocalMux I__5194 (
            .O(N__29879),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__5193 (
            .O(N__29874),
            .I(N__29868));
    InMux I__5192 (
            .O(N__29873),
            .I(N__29868));
    LocalMux I__5191 (
            .O(N__29868),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    InMux I__5190 (
            .O(N__29865),
            .I(N__29862));
    LocalMux I__5189 (
            .O(N__29862),
            .I(N__29858));
    InMux I__5188 (
            .O(N__29861),
            .I(N__29855));
    Span4Mux_v I__5187 (
            .O(N__29858),
            .I(N__29852));
    LocalMux I__5186 (
            .O(N__29855),
            .I(N__29849));
    Sp12to4 I__5185 (
            .O(N__29852),
            .I(N__29844));
    Span12Mux_v I__5184 (
            .O(N__29849),
            .I(N__29844));
    Odrv12 I__5183 (
            .O(N__29844),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    InMux I__5182 (
            .O(N__29841),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ));
    InMux I__5181 (
            .O(N__29838),
            .I(N__29835));
    LocalMux I__5180 (
            .O(N__29835),
            .I(N__29831));
    InMux I__5179 (
            .O(N__29834),
            .I(N__29828));
    Span4Mux_s2_h I__5178 (
            .O(N__29831),
            .I(N__29825));
    LocalMux I__5177 (
            .O(N__29828),
            .I(N__29822));
    Span4Mux_v I__5176 (
            .O(N__29825),
            .I(N__29819));
    Span4Mux_v I__5175 (
            .O(N__29822),
            .I(N__29814));
    Span4Mux_h I__5174 (
            .O(N__29819),
            .I(N__29814));
    Odrv4 I__5173 (
            .O(N__29814),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    InMux I__5172 (
            .O(N__29811),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ));
    InMux I__5171 (
            .O(N__29808),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ));
    InMux I__5170 (
            .O(N__29805),
            .I(N__29802));
    LocalMux I__5169 (
            .O(N__29802),
            .I(N__29799));
    Odrv12 I__5168 (
            .O(N__29799),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_31 ));
    InMux I__5167 (
            .O(N__29796),
            .I(N__29793));
    LocalMux I__5166 (
            .O(N__29793),
            .I(N__29790));
    Odrv12 I__5165 (
            .O(N__29790),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ));
    InMux I__5164 (
            .O(N__29787),
            .I(N__29779));
    InMux I__5163 (
            .O(N__29786),
            .I(N__29768));
    InMux I__5162 (
            .O(N__29785),
            .I(N__29768));
    InMux I__5161 (
            .O(N__29784),
            .I(N__29768));
    InMux I__5160 (
            .O(N__29783),
            .I(N__29768));
    InMux I__5159 (
            .O(N__29782),
            .I(N__29768));
    LocalMux I__5158 (
            .O(N__29779),
            .I(N__29765));
    LocalMux I__5157 (
            .O(N__29768),
            .I(N__29759));
    Span4Mux_h I__5156 (
            .O(N__29765),
            .I(N__29755));
    InMux I__5155 (
            .O(N__29764),
            .I(N__29748));
    InMux I__5154 (
            .O(N__29763),
            .I(N__29748));
    InMux I__5153 (
            .O(N__29762),
            .I(N__29748));
    Span4Mux_s3_h I__5152 (
            .O(N__29759),
            .I(N__29745));
    InMux I__5151 (
            .O(N__29758),
            .I(N__29742));
    Span4Mux_h I__5150 (
            .O(N__29755),
            .I(N__29737));
    LocalMux I__5149 (
            .O(N__29748),
            .I(N__29737));
    Odrv4 I__5148 (
            .O(N__29745),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    LocalMux I__5147 (
            .O(N__29742),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__5146 (
            .O(N__29737),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__5145 (
            .O(N__29730),
            .I(N__29727));
    LocalMux I__5144 (
            .O(N__29727),
            .I(N__29724));
    Odrv12 I__5143 (
            .O(N__29724),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__5142 (
            .O(N__29721),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__5141 (
            .O(N__29718),
            .I(N__29715));
    LocalMux I__5140 (
            .O(N__29715),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    InMux I__5139 (
            .O(N__29712),
            .I(N__29708));
    InMux I__5138 (
            .O(N__29711),
            .I(N__29705));
    LocalMux I__5137 (
            .O(N__29708),
            .I(N__29702));
    LocalMux I__5136 (
            .O(N__29705),
            .I(N__29699));
    Span12Mux_s9_h I__5135 (
            .O(N__29702),
            .I(N__29696));
    Span12Mux_v I__5134 (
            .O(N__29699),
            .I(N__29693));
    Odrv12 I__5133 (
            .O(N__29696),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    Odrv12 I__5132 (
            .O(N__29693),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__5131 (
            .O(N__29688),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__5130 (
            .O(N__29685),
            .I(N__29682));
    LocalMux I__5129 (
            .O(N__29682),
            .I(N__29679));
    Span4Mux_s2_h I__5128 (
            .O(N__29679),
            .I(N__29675));
    InMux I__5127 (
            .O(N__29678),
            .I(N__29672));
    Span4Mux_h I__5126 (
            .O(N__29675),
            .I(N__29669));
    LocalMux I__5125 (
            .O(N__29672),
            .I(N__29666));
    Span4Mux_h I__5124 (
            .O(N__29669),
            .I(N__29663));
    Odrv12 I__5123 (
            .O(N__29666),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    Odrv4 I__5122 (
            .O(N__29663),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    InMux I__5121 (
            .O(N__29658),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    InMux I__5120 (
            .O(N__29655),
            .I(N__29651));
    InMux I__5119 (
            .O(N__29654),
            .I(N__29648));
    LocalMux I__5118 (
            .O(N__29651),
            .I(N__29645));
    LocalMux I__5117 (
            .O(N__29648),
            .I(N__29642));
    Span4Mux_v I__5116 (
            .O(N__29645),
            .I(N__29637));
    Span4Mux_v I__5115 (
            .O(N__29642),
            .I(N__29637));
    Sp12to4 I__5114 (
            .O(N__29637),
            .I(N__29634));
    Odrv12 I__5113 (
            .O(N__29634),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__5112 (
            .O(N__29631),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__5111 (
            .O(N__29628),
            .I(N__29625));
    LocalMux I__5110 (
            .O(N__29625),
            .I(N__29621));
    InMux I__5109 (
            .O(N__29624),
            .I(N__29618));
    Span4Mux_h I__5108 (
            .O(N__29621),
            .I(N__29615));
    LocalMux I__5107 (
            .O(N__29618),
            .I(N__29612));
    Span4Mux_h I__5106 (
            .O(N__29615),
            .I(N__29609));
    Span12Mux_s9_h I__5105 (
            .O(N__29612),
            .I(N__29606));
    Odrv4 I__5104 (
            .O(N__29609),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    Odrv12 I__5103 (
            .O(N__29606),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__5102 (
            .O(N__29601),
            .I(bfn_9_16_0_));
    InMux I__5101 (
            .O(N__29598),
            .I(N__29595));
    LocalMux I__5100 (
            .O(N__29595),
            .I(N__29591));
    InMux I__5099 (
            .O(N__29594),
            .I(N__29588));
    Span4Mux_s1_h I__5098 (
            .O(N__29591),
            .I(N__29585));
    LocalMux I__5097 (
            .O(N__29588),
            .I(N__29582));
    Span4Mux_h I__5096 (
            .O(N__29585),
            .I(N__29579));
    Span12Mux_v I__5095 (
            .O(N__29582),
            .I(N__29576));
    Span4Mux_h I__5094 (
            .O(N__29579),
            .I(N__29573));
    Odrv12 I__5093 (
            .O(N__29576),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    Odrv4 I__5092 (
            .O(N__29573),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__5091 (
            .O(N__29568),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__5090 (
            .O(N__29565),
            .I(N__29561));
    InMux I__5089 (
            .O(N__29564),
            .I(N__29558));
    LocalMux I__5088 (
            .O(N__29561),
            .I(N__29555));
    LocalMux I__5087 (
            .O(N__29558),
            .I(N__29552));
    Span4Mux_s1_h I__5086 (
            .O(N__29555),
            .I(N__29549));
    Span4Mux_v I__5085 (
            .O(N__29552),
            .I(N__29546));
    Span4Mux_h I__5084 (
            .O(N__29549),
            .I(N__29543));
    Span4Mux_h I__5083 (
            .O(N__29546),
            .I(N__29538));
    Span4Mux_h I__5082 (
            .O(N__29543),
            .I(N__29538));
    Odrv4 I__5081 (
            .O(N__29538),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__5080 (
            .O(N__29535),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__5079 (
            .O(N__29532),
            .I(N__29528));
    InMux I__5078 (
            .O(N__29531),
            .I(N__29525));
    LocalMux I__5077 (
            .O(N__29528),
            .I(N__29522));
    LocalMux I__5076 (
            .O(N__29525),
            .I(N__29519));
    Span4Mux_s1_h I__5075 (
            .O(N__29522),
            .I(N__29516));
    Span4Mux_v I__5074 (
            .O(N__29519),
            .I(N__29513));
    Span4Mux_h I__5073 (
            .O(N__29516),
            .I(N__29510));
    Span4Mux_h I__5072 (
            .O(N__29513),
            .I(N__29505));
    Span4Mux_h I__5071 (
            .O(N__29510),
            .I(N__29505));
    Odrv4 I__5070 (
            .O(N__29505),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    InMux I__5069 (
            .O(N__29502),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ));
    InMux I__5068 (
            .O(N__29499),
            .I(N__29496));
    LocalMux I__5067 (
            .O(N__29496),
            .I(N__29493));
    Span4Mux_s1_h I__5066 (
            .O(N__29493),
            .I(N__29489));
    InMux I__5065 (
            .O(N__29492),
            .I(N__29486));
    Span4Mux_h I__5064 (
            .O(N__29489),
            .I(N__29483));
    LocalMux I__5063 (
            .O(N__29486),
            .I(N__29480));
    Span4Mux_h I__5062 (
            .O(N__29483),
            .I(N__29477));
    Odrv12 I__5061 (
            .O(N__29480),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    Odrv4 I__5060 (
            .O(N__29477),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    InMux I__5059 (
            .O(N__29472),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ));
    InMux I__5058 (
            .O(N__29469),
            .I(N__29465));
    InMux I__5057 (
            .O(N__29468),
            .I(N__29462));
    LocalMux I__5056 (
            .O(N__29465),
            .I(N__29459));
    LocalMux I__5055 (
            .O(N__29462),
            .I(N__29456));
    Span12Mux_s9_h I__5054 (
            .O(N__29459),
            .I(N__29453));
    Odrv12 I__5053 (
            .O(N__29456),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv12 I__5052 (
            .O(N__29453),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__5051 (
            .O(N__29448),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__5050 (
            .O(N__29445),
            .I(N__29441));
    InMux I__5049 (
            .O(N__29444),
            .I(N__29438));
    LocalMux I__5048 (
            .O(N__29441),
            .I(N__29435));
    LocalMux I__5047 (
            .O(N__29438),
            .I(N__29432));
    Span4Mux_v I__5046 (
            .O(N__29435),
            .I(N__29429));
    Span4Mux_v I__5045 (
            .O(N__29432),
            .I(N__29424));
    Span4Mux_v I__5044 (
            .O(N__29429),
            .I(N__29424));
    Sp12to4 I__5043 (
            .O(N__29424),
            .I(N__29421));
    Odrv12 I__5042 (
            .O(N__29421),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__5041 (
            .O(N__29418),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__5040 (
            .O(N__29415),
            .I(N__29412));
    LocalMux I__5039 (
            .O(N__29412),
            .I(N__29408));
    InMux I__5038 (
            .O(N__29411),
            .I(N__29405));
    Span4Mux_v I__5037 (
            .O(N__29408),
            .I(N__29402));
    LocalMux I__5036 (
            .O(N__29405),
            .I(N__29397));
    Sp12to4 I__5035 (
            .O(N__29402),
            .I(N__29397));
    Odrv12 I__5034 (
            .O(N__29397),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__5033 (
            .O(N__29394),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__5032 (
            .O(N__29391),
            .I(N__29387));
    InMux I__5031 (
            .O(N__29390),
            .I(N__29384));
    LocalMux I__5030 (
            .O(N__29387),
            .I(N__29381));
    LocalMux I__5029 (
            .O(N__29384),
            .I(N__29378));
    Span4Mux_s1_h I__5028 (
            .O(N__29381),
            .I(N__29375));
    Span4Mux_v I__5027 (
            .O(N__29378),
            .I(N__29372));
    Span4Mux_h I__5026 (
            .O(N__29375),
            .I(N__29369));
    Span4Mux_h I__5025 (
            .O(N__29372),
            .I(N__29364));
    Span4Mux_h I__5024 (
            .O(N__29369),
            .I(N__29364));
    Odrv4 I__5023 (
            .O(N__29364),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__5022 (
            .O(N__29361),
            .I(bfn_9_15_0_));
    InMux I__5021 (
            .O(N__29358),
            .I(N__29354));
    InMux I__5020 (
            .O(N__29357),
            .I(N__29351));
    LocalMux I__5019 (
            .O(N__29354),
            .I(N__29348));
    LocalMux I__5018 (
            .O(N__29351),
            .I(N__29345));
    Span12Mux_s9_h I__5017 (
            .O(N__29348),
            .I(N__29342));
    Odrv12 I__5016 (
            .O(N__29345),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    Odrv12 I__5015 (
            .O(N__29342),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__5014 (
            .O(N__29337),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__5013 (
            .O(N__29334),
            .I(N__29331));
    LocalMux I__5012 (
            .O(N__29331),
            .I(N__29328));
    Span4Mux_s1_h I__5011 (
            .O(N__29328),
            .I(N__29324));
    InMux I__5010 (
            .O(N__29327),
            .I(N__29321));
    Span4Mux_h I__5009 (
            .O(N__29324),
            .I(N__29318));
    LocalMux I__5008 (
            .O(N__29321),
            .I(N__29315));
    Span4Mux_h I__5007 (
            .O(N__29318),
            .I(N__29312));
    Odrv12 I__5006 (
            .O(N__29315),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    Odrv4 I__5005 (
            .O(N__29312),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__5004 (
            .O(N__29307),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__5003 (
            .O(N__29304),
            .I(N__29300));
    InMux I__5002 (
            .O(N__29303),
            .I(N__29297));
    LocalMux I__5001 (
            .O(N__29300),
            .I(N__29294));
    LocalMux I__5000 (
            .O(N__29297),
            .I(N__29291));
    Span4Mux_s1_h I__4999 (
            .O(N__29294),
            .I(N__29288));
    Span4Mux_v I__4998 (
            .O(N__29291),
            .I(N__29285));
    Span4Mux_h I__4997 (
            .O(N__29288),
            .I(N__29282));
    Span4Mux_h I__4996 (
            .O(N__29285),
            .I(N__29277));
    Span4Mux_h I__4995 (
            .O(N__29282),
            .I(N__29277));
    Odrv4 I__4994 (
            .O(N__29277),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    InMux I__4993 (
            .O(N__29274),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__4992 (
            .O(N__29271),
            .I(N__29267));
    InMux I__4991 (
            .O(N__29270),
            .I(N__29264));
    LocalMux I__4990 (
            .O(N__29267),
            .I(N__29261));
    LocalMux I__4989 (
            .O(N__29264),
            .I(N__29258));
    Span4Mux_v I__4988 (
            .O(N__29261),
            .I(N__29253));
    Span4Mux_v I__4987 (
            .O(N__29258),
            .I(N__29253));
    Sp12to4 I__4986 (
            .O(N__29253),
            .I(N__29250));
    Odrv12 I__4985 (
            .O(N__29250),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    InMux I__4984 (
            .O(N__29247),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__4983 (
            .O(N__29244),
            .I(N__29240));
    InMux I__4982 (
            .O(N__29243),
            .I(N__29237));
    LocalMux I__4981 (
            .O(N__29240),
            .I(N__29234));
    LocalMux I__4980 (
            .O(N__29237),
            .I(N__29231));
    Span4Mux_v I__4979 (
            .O(N__29234),
            .I(N__29228));
    Sp12to4 I__4978 (
            .O(N__29231),
            .I(N__29225));
    Sp12to4 I__4977 (
            .O(N__29228),
            .I(N__29220));
    Span12Mux_v I__4976 (
            .O(N__29225),
            .I(N__29220));
    Odrv12 I__4975 (
            .O(N__29220),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__4974 (
            .O(N__29217),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__4973 (
            .O(N__29214),
            .I(N__29210));
    InMux I__4972 (
            .O(N__29213),
            .I(N__29207));
    LocalMux I__4971 (
            .O(N__29210),
            .I(N__29204));
    LocalMux I__4970 (
            .O(N__29207),
            .I(N__29199));
    Span12Mux_v I__4969 (
            .O(N__29204),
            .I(N__29199));
    Odrv12 I__4968 (
            .O(N__29199),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__4967 (
            .O(N__29196),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__4966 (
            .O(N__29193),
            .I(N__29189));
    InMux I__4965 (
            .O(N__29192),
            .I(N__29186));
    LocalMux I__4964 (
            .O(N__29189),
            .I(N__29183));
    LocalMux I__4963 (
            .O(N__29186),
            .I(N__29180));
    Span12Mux_s9_h I__4962 (
            .O(N__29183),
            .I(N__29177));
    Odrv12 I__4961 (
            .O(N__29180),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv12 I__4960 (
            .O(N__29177),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__4959 (
            .O(N__29172),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__4958 (
            .O(N__29169),
            .I(N__29166));
    LocalMux I__4957 (
            .O(N__29166),
            .I(N__29163));
    Span4Mux_v I__4956 (
            .O(N__29163),
            .I(N__29159));
    InMux I__4955 (
            .O(N__29162),
            .I(N__29156));
    Span4Mux_h I__4954 (
            .O(N__29159),
            .I(N__29153));
    LocalMux I__4953 (
            .O(N__29156),
            .I(N__29150));
    Span4Mux_h I__4952 (
            .O(N__29153),
            .I(N__29147));
    Odrv12 I__4951 (
            .O(N__29150),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__4950 (
            .O(N__29147),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__4949 (
            .O(N__29142),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__4948 (
            .O(N__29139),
            .I(N__29136));
    LocalMux I__4947 (
            .O(N__29136),
            .I(N__29132));
    InMux I__4946 (
            .O(N__29135),
            .I(N__29129));
    Span4Mux_v I__4945 (
            .O(N__29132),
            .I(N__29126));
    LocalMux I__4944 (
            .O(N__29129),
            .I(N__29123));
    Sp12to4 I__4943 (
            .O(N__29126),
            .I(N__29120));
    Span4Mux_h I__4942 (
            .O(N__29123),
            .I(N__29117));
    Span12Mux_s9_h I__4941 (
            .O(N__29120),
            .I(N__29114));
    Odrv4 I__4940 (
            .O(N__29117),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv12 I__4939 (
            .O(N__29114),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__4938 (
            .O(N__29109),
            .I(bfn_9_14_0_));
    InMux I__4937 (
            .O(N__29106),
            .I(N__29103));
    LocalMux I__4936 (
            .O(N__29103),
            .I(N__29099));
    InMux I__4935 (
            .O(N__29102),
            .I(N__29096));
    Span4Mux_h I__4934 (
            .O(N__29099),
            .I(N__29093));
    LocalMux I__4933 (
            .O(N__29096),
            .I(N__29090));
    Sp12to4 I__4932 (
            .O(N__29093),
            .I(N__29087));
    Span12Mux_s4_h I__4931 (
            .O(N__29090),
            .I(N__29082));
    Span12Mux_v I__4930 (
            .O(N__29087),
            .I(N__29082));
    Odrv12 I__4929 (
            .O(N__29082),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__4928 (
            .O(N__29079),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__4927 (
            .O(N__29076),
            .I(N__29073));
    LocalMux I__4926 (
            .O(N__29073),
            .I(N__29069));
    InMux I__4925 (
            .O(N__29072),
            .I(N__29066));
    Span4Mux_v I__4924 (
            .O(N__29069),
            .I(N__29063));
    LocalMux I__4923 (
            .O(N__29066),
            .I(N__29060));
    Span4Mux_h I__4922 (
            .O(N__29063),
            .I(N__29057));
    Span12Mux_v I__4921 (
            .O(N__29060),
            .I(N__29054));
    Span4Mux_h I__4920 (
            .O(N__29057),
            .I(N__29051));
    Odrv12 I__4919 (
            .O(N__29054),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__4918 (
            .O(N__29051),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__4917 (
            .O(N__29046),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__4916 (
            .O(N__29043),
            .I(N__29040));
    LocalMux I__4915 (
            .O(N__29040),
            .I(N__29036));
    InMux I__4914 (
            .O(N__29039),
            .I(N__29033));
    Span4Mux_v I__4913 (
            .O(N__29036),
            .I(N__29030));
    LocalMux I__4912 (
            .O(N__29033),
            .I(N__29027));
    Span4Mux_h I__4911 (
            .O(N__29030),
            .I(N__29024));
    Span12Mux_s9_h I__4910 (
            .O(N__29027),
            .I(N__29021));
    Span4Mux_h I__4909 (
            .O(N__29024),
            .I(N__29018));
    Odrv12 I__4908 (
            .O(N__29021),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__4907 (
            .O(N__29018),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__4906 (
            .O(N__29013),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__4905 (
            .O(N__29010),
            .I(N__29006));
    InMux I__4904 (
            .O(N__29009),
            .I(N__29003));
    LocalMux I__4903 (
            .O(N__29006),
            .I(N__29000));
    LocalMux I__4902 (
            .O(N__29003),
            .I(N__28997));
    Span4Mux_v I__4901 (
            .O(N__29000),
            .I(N__28994));
    Span4Mux_v I__4900 (
            .O(N__28997),
            .I(N__28991));
    Span4Mux_h I__4899 (
            .O(N__28994),
            .I(N__28988));
    Span4Mux_h I__4898 (
            .O(N__28991),
            .I(N__28985));
    Span4Mux_h I__4897 (
            .O(N__28988),
            .I(N__28982));
    Odrv4 I__4896 (
            .O(N__28985),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__4895 (
            .O(N__28982),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__4894 (
            .O(N__28977),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__4893 (
            .O(N__28974),
            .I(N__28970));
    InMux I__4892 (
            .O(N__28973),
            .I(N__28967));
    LocalMux I__4891 (
            .O(N__28970),
            .I(N__28962));
    LocalMux I__4890 (
            .O(N__28967),
            .I(N__28959));
    InMux I__4889 (
            .O(N__28966),
            .I(N__28954));
    InMux I__4888 (
            .O(N__28965),
            .I(N__28954));
    Span4Mux_v I__4887 (
            .O(N__28962),
            .I(N__28951));
    Span4Mux_h I__4886 (
            .O(N__28959),
            .I(N__28948));
    LocalMux I__4885 (
            .O(N__28954),
            .I(N__28945));
    Odrv4 I__4884 (
            .O(N__28951),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__4883 (
            .O(N__28948),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv12 I__4882 (
            .O(N__28945),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__4881 (
            .O(N__28938),
            .I(N__28933));
    InMux I__4880 (
            .O(N__28937),
            .I(N__28930));
    InMux I__4879 (
            .O(N__28936),
            .I(N__28927));
    LocalMux I__4878 (
            .O(N__28933),
            .I(N__28924));
    LocalMux I__4877 (
            .O(N__28930),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__4876 (
            .O(N__28927),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__4875 (
            .O(N__28924),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__4874 (
            .O(N__28917),
            .I(N__28911));
    InMux I__4873 (
            .O(N__28916),
            .I(N__28911));
    LocalMux I__4872 (
            .O(N__28911),
            .I(N__28906));
    InMux I__4871 (
            .O(N__28910),
            .I(N__28903));
    InMux I__4870 (
            .O(N__28909),
            .I(N__28900));
    Span4Mux_h I__4869 (
            .O(N__28906),
            .I(N__28897));
    LocalMux I__4868 (
            .O(N__28903),
            .I(N__28894));
    LocalMux I__4867 (
            .O(N__28900),
            .I(N__28887));
    Span4Mux_v I__4866 (
            .O(N__28897),
            .I(N__28887));
    Span4Mux_h I__4865 (
            .O(N__28894),
            .I(N__28887));
    Odrv4 I__4864 (
            .O(N__28887),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__4863 (
            .O(N__28884),
            .I(N__28881));
    LocalMux I__4862 (
            .O(N__28881),
            .I(N__28878));
    Span4Mux_v I__4861 (
            .O(N__28878),
            .I(N__28874));
    InMux I__4860 (
            .O(N__28877),
            .I(N__28871));
    Odrv4 I__4859 (
            .O(N__28874),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    LocalMux I__4858 (
            .O(N__28871),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    InMux I__4857 (
            .O(N__28866),
            .I(N__28861));
    InMux I__4856 (
            .O(N__28865),
            .I(N__28858));
    InMux I__4855 (
            .O(N__28864),
            .I(N__28855));
    LocalMux I__4854 (
            .O(N__28861),
            .I(N__28852));
    LocalMux I__4853 (
            .O(N__28858),
            .I(N__28849));
    LocalMux I__4852 (
            .O(N__28855),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv4 I__4851 (
            .O(N__28852),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv4 I__4850 (
            .O(N__28849),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    InMux I__4849 (
            .O(N__28842),
            .I(N__28835));
    InMux I__4848 (
            .O(N__28841),
            .I(N__28835));
    InMux I__4847 (
            .O(N__28840),
            .I(N__28831));
    LocalMux I__4846 (
            .O(N__28835),
            .I(N__28828));
    InMux I__4845 (
            .O(N__28834),
            .I(N__28825));
    LocalMux I__4844 (
            .O(N__28831),
            .I(N__28820));
    Span4Mux_v I__4843 (
            .O(N__28828),
            .I(N__28820));
    LocalMux I__4842 (
            .O(N__28825),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv4 I__4841 (
            .O(N__28820),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    CascadeMux I__4840 (
            .O(N__28815),
            .I(N__28812));
    InMux I__4839 (
            .O(N__28812),
            .I(N__28806));
    InMux I__4838 (
            .O(N__28811),
            .I(N__28806));
    LocalMux I__4837 (
            .O(N__28806),
            .I(N__28803));
    Odrv4 I__4836 (
            .O(N__28803),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    InMux I__4835 (
            .O(N__28800),
            .I(N__28795));
    InMux I__4834 (
            .O(N__28799),
            .I(N__28792));
    InMux I__4833 (
            .O(N__28798),
            .I(N__28789));
    LocalMux I__4832 (
            .O(N__28795),
            .I(N__28786));
    LocalMux I__4831 (
            .O(N__28792),
            .I(N__28783));
    LocalMux I__4830 (
            .O(N__28789),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__4829 (
            .O(N__28786),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__4828 (
            .O(N__28783),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    InMux I__4827 (
            .O(N__28776),
            .I(N__28772));
    CascadeMux I__4826 (
            .O(N__28775),
            .I(N__28769));
    LocalMux I__4825 (
            .O(N__28772),
            .I(N__28765));
    InMux I__4824 (
            .O(N__28769),
            .I(N__28762));
    InMux I__4823 (
            .O(N__28768),
            .I(N__28759));
    Span4Mux_h I__4822 (
            .O(N__28765),
            .I(N__28751));
    LocalMux I__4821 (
            .O(N__28762),
            .I(N__28751));
    LocalMux I__4820 (
            .O(N__28759),
            .I(N__28751));
    InMux I__4819 (
            .O(N__28758),
            .I(N__28748));
    Span4Mux_v I__4818 (
            .O(N__28751),
            .I(N__28745));
    LocalMux I__4817 (
            .O(N__28748),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__4816 (
            .O(N__28745),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__4815 (
            .O(N__28740),
            .I(N__28737));
    LocalMux I__4814 (
            .O(N__28737),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__4813 (
            .O(N__28734),
            .I(N__28730));
    InMux I__4812 (
            .O(N__28733),
            .I(N__28727));
    LocalMux I__4811 (
            .O(N__28730),
            .I(N__28724));
    LocalMux I__4810 (
            .O(N__28727),
            .I(N__28721));
    Span4Mux_h I__4809 (
            .O(N__28724),
            .I(N__28718));
    Span4Mux_v I__4808 (
            .O(N__28721),
            .I(N__28715));
    Span4Mux_h I__4807 (
            .O(N__28718),
            .I(N__28712));
    Span4Mux_h I__4806 (
            .O(N__28715),
            .I(N__28709));
    Span4Mux_v I__4805 (
            .O(N__28712),
            .I(N__28706));
    Span4Mux_h I__4804 (
            .O(N__28709),
            .I(N__28703));
    Odrv4 I__4803 (
            .O(N__28706),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    Odrv4 I__4802 (
            .O(N__28703),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__4801 (
            .O(N__28698),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__4800 (
            .O(N__28695),
            .I(N__28692));
    LocalMux I__4799 (
            .O(N__28692),
            .I(N__28689));
    Span4Mux_v I__4798 (
            .O(N__28689),
            .I(N__28685));
    InMux I__4797 (
            .O(N__28688),
            .I(N__28682));
    Span4Mux_h I__4796 (
            .O(N__28685),
            .I(N__28679));
    LocalMux I__4795 (
            .O(N__28682),
            .I(N__28676));
    Span4Mux_h I__4794 (
            .O(N__28679),
            .I(N__28673));
    Odrv12 I__4793 (
            .O(N__28676),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv4 I__4792 (
            .O(N__28673),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__4791 (
            .O(N__28668),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__4790 (
            .O(N__28665),
            .I(N__28661));
    InMux I__4789 (
            .O(N__28664),
            .I(N__28658));
    LocalMux I__4788 (
            .O(N__28661),
            .I(N__28655));
    LocalMux I__4787 (
            .O(N__28658),
            .I(N__28652));
    Span4Mux_v I__4786 (
            .O(N__28655),
            .I(N__28649));
    Span4Mux_h I__4785 (
            .O(N__28652),
            .I(N__28646));
    Span4Mux_h I__4784 (
            .O(N__28649),
            .I(N__28643));
    Span4Mux_h I__4783 (
            .O(N__28646),
            .I(N__28638));
    Span4Mux_h I__4782 (
            .O(N__28643),
            .I(N__28638));
    Odrv4 I__4781 (
            .O(N__28638),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__4780 (
            .O(N__28635),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__4779 (
            .O(N__28632),
            .I(N__28628));
    InMux I__4778 (
            .O(N__28631),
            .I(N__28624));
    LocalMux I__4777 (
            .O(N__28628),
            .I(N__28621));
    InMux I__4776 (
            .O(N__28627),
            .I(N__28618));
    LocalMux I__4775 (
            .O(N__28624),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    Odrv12 I__4774 (
            .O(N__28621),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    LocalMux I__4773 (
            .O(N__28618),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__4772 (
            .O(N__28611),
            .I(N__28606));
    CascadeMux I__4771 (
            .O(N__28610),
            .I(N__28602));
    InMux I__4770 (
            .O(N__28609),
            .I(N__28599));
    LocalMux I__4769 (
            .O(N__28606),
            .I(N__28596));
    InMux I__4768 (
            .O(N__28605),
            .I(N__28593));
    InMux I__4767 (
            .O(N__28602),
            .I(N__28590));
    LocalMux I__4766 (
            .O(N__28599),
            .I(N__28587));
    Span4Mux_h I__4765 (
            .O(N__28596),
            .I(N__28580));
    LocalMux I__4764 (
            .O(N__28593),
            .I(N__28580));
    LocalMux I__4763 (
            .O(N__28590),
            .I(N__28580));
    Span4Mux_h I__4762 (
            .O(N__28587),
            .I(N__28575));
    Span4Mux_v I__4761 (
            .O(N__28580),
            .I(N__28575));
    Odrv4 I__4760 (
            .O(N__28575),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__4759 (
            .O(N__28572),
            .I(N__28566));
    InMux I__4758 (
            .O(N__28571),
            .I(N__28566));
    LocalMux I__4757 (
            .O(N__28566),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    InMux I__4756 (
            .O(N__28563),
            .I(N__28559));
    InMux I__4755 (
            .O(N__28562),
            .I(N__28555));
    LocalMux I__4754 (
            .O(N__28559),
            .I(N__28552));
    InMux I__4753 (
            .O(N__28558),
            .I(N__28549));
    LocalMux I__4752 (
            .O(N__28555),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    Odrv4 I__4751 (
            .O(N__28552),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__4750 (
            .O(N__28549),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    CascadeMux I__4749 (
            .O(N__28542),
            .I(N__28537));
    InMux I__4748 (
            .O(N__28541),
            .I(N__28533));
    InMux I__4747 (
            .O(N__28540),
            .I(N__28528));
    InMux I__4746 (
            .O(N__28537),
            .I(N__28528));
    InMux I__4745 (
            .O(N__28536),
            .I(N__28525));
    LocalMux I__4744 (
            .O(N__28533),
            .I(N__28520));
    LocalMux I__4743 (
            .O(N__28528),
            .I(N__28520));
    LocalMux I__4742 (
            .O(N__28525),
            .I(N__28517));
    Span4Mux_v I__4741 (
            .O(N__28520),
            .I(N__28514));
    Odrv4 I__4740 (
            .O(N__28517),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__4739 (
            .O(N__28514),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__4738 (
            .O(N__28509),
            .I(N__28505));
    InMux I__4737 (
            .O(N__28508),
            .I(N__28501));
    LocalMux I__4736 (
            .O(N__28505),
            .I(N__28498));
    InMux I__4735 (
            .O(N__28504),
            .I(N__28495));
    LocalMux I__4734 (
            .O(N__28501),
            .I(N__28492));
    Span4Mux_h I__4733 (
            .O(N__28498),
            .I(N__28489));
    LocalMux I__4732 (
            .O(N__28495),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv12 I__4731 (
            .O(N__28492),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv4 I__4730 (
            .O(N__28489),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__4729 (
            .O(N__28482),
            .I(N__28478));
    InMux I__4728 (
            .O(N__28481),
            .I(N__28474));
    LocalMux I__4727 (
            .O(N__28478),
            .I(N__28471));
    CascadeMux I__4726 (
            .O(N__28477),
            .I(N__28467));
    LocalMux I__4725 (
            .O(N__28474),
            .I(N__28464));
    Span4Mux_h I__4724 (
            .O(N__28471),
            .I(N__28461));
    InMux I__4723 (
            .O(N__28470),
            .I(N__28458));
    InMux I__4722 (
            .O(N__28467),
            .I(N__28455));
    Odrv12 I__4721 (
            .O(N__28464),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv4 I__4720 (
            .O(N__28461),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__4719 (
            .O(N__28458),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__4718 (
            .O(N__28455),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__4717 (
            .O(N__28446),
            .I(N__28440));
    InMux I__4716 (
            .O(N__28445),
            .I(N__28440));
    LocalMux I__4715 (
            .O(N__28440),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    InMux I__4714 (
            .O(N__28437),
            .I(N__28434));
    LocalMux I__4713 (
            .O(N__28434),
            .I(N__28431));
    Span4Mux_s1_v I__4712 (
            .O(N__28431),
            .I(N__28427));
    InMux I__4711 (
            .O(N__28430),
            .I(N__28424));
    Span4Mux_v I__4710 (
            .O(N__28427),
            .I(N__28419));
    LocalMux I__4709 (
            .O(N__28424),
            .I(N__28416));
    InMux I__4708 (
            .O(N__28423),
            .I(N__28413));
    InMux I__4707 (
            .O(N__28422),
            .I(N__28410));
    Span4Mux_v I__4706 (
            .O(N__28419),
            .I(N__28407));
    Span4Mux_h I__4705 (
            .O(N__28416),
            .I(N__28402));
    LocalMux I__4704 (
            .O(N__28413),
            .I(N__28402));
    LocalMux I__4703 (
            .O(N__28410),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__4702 (
            .O(N__28407),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__4701 (
            .O(N__28402),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__4700 (
            .O(N__28395),
            .I(N__28390));
    InMux I__4699 (
            .O(N__28394),
            .I(N__28387));
    InMux I__4698 (
            .O(N__28393),
            .I(N__28384));
    LocalMux I__4697 (
            .O(N__28390),
            .I(N__28381));
    LocalMux I__4696 (
            .O(N__28387),
            .I(N__28378));
    LocalMux I__4695 (
            .O(N__28384),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    Odrv12 I__4694 (
            .O(N__28381),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    Odrv4 I__4693 (
            .O(N__28378),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    InMux I__4692 (
            .O(N__28371),
            .I(N__28368));
    LocalMux I__4691 (
            .O(N__28368),
            .I(N__28365));
    Span4Mux_v I__4690 (
            .O(N__28365),
            .I(N__28359));
    InMux I__4689 (
            .O(N__28364),
            .I(N__28356));
    InMux I__4688 (
            .O(N__28363),
            .I(N__28351));
    InMux I__4687 (
            .O(N__28362),
            .I(N__28351));
    Odrv4 I__4686 (
            .O(N__28359),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__4685 (
            .O(N__28356),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__4684 (
            .O(N__28351),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__4683 (
            .O(N__28344),
            .I(N__28340));
    InMux I__4682 (
            .O(N__28343),
            .I(N__28336));
    LocalMux I__4681 (
            .O(N__28340),
            .I(N__28333));
    InMux I__4680 (
            .O(N__28339),
            .I(N__28330));
    LocalMux I__4679 (
            .O(N__28336),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv12 I__4678 (
            .O(N__28333),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    LocalMux I__4677 (
            .O(N__28330),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    CascadeMux I__4676 (
            .O(N__28323),
            .I(N__28320));
    InMux I__4675 (
            .O(N__28320),
            .I(N__28314));
    InMux I__4674 (
            .O(N__28319),
            .I(N__28314));
    LocalMux I__4673 (
            .O(N__28314),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    InMux I__4672 (
            .O(N__28311),
            .I(N__28308));
    LocalMux I__4671 (
            .O(N__28308),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    InMux I__4670 (
            .O(N__28305),
            .I(N__28302));
    LocalMux I__4669 (
            .O(N__28302),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    CascadeMux I__4668 (
            .O(N__28299),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_ ));
    InMux I__4667 (
            .O(N__28296),
            .I(N__28293));
    LocalMux I__4666 (
            .O(N__28293),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__4665 (
            .O(N__28290),
            .I(N__28287));
    LocalMux I__4664 (
            .O(N__28287),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    CascadeMux I__4663 (
            .O(N__28284),
            .I(N__28281));
    InMux I__4662 (
            .O(N__28281),
            .I(N__28275));
    InMux I__4661 (
            .O(N__28280),
            .I(N__28275));
    LocalMux I__4660 (
            .O(N__28275),
            .I(N__28272));
    Odrv4 I__4659 (
            .O(N__28272),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    CascadeMux I__4658 (
            .O(N__28269),
            .I(N__28266));
    InMux I__4657 (
            .O(N__28266),
            .I(N__28259));
    InMux I__4656 (
            .O(N__28265),
            .I(N__28259));
    InMux I__4655 (
            .O(N__28264),
            .I(N__28256));
    LocalMux I__4654 (
            .O(N__28259),
            .I(N__28253));
    LocalMux I__4653 (
            .O(N__28256),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__4652 (
            .O(N__28253),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__4651 (
            .O(N__28248),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__4650 (
            .O(N__28245),
            .I(N__28240));
    InMux I__4649 (
            .O(N__28244),
            .I(N__28235));
    InMux I__4648 (
            .O(N__28243),
            .I(N__28235));
    LocalMux I__4647 (
            .O(N__28240),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__4646 (
            .O(N__28235),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__4645 (
            .O(N__28230),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__4644 (
            .O(N__28227),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__4643 (
            .O(N__28224),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__4642 (
            .O(N__28221),
            .I(N__28217));
    InMux I__4641 (
            .O(N__28220),
            .I(N__28213));
    LocalMux I__4640 (
            .O(N__28217),
            .I(N__28210));
    InMux I__4639 (
            .O(N__28216),
            .I(N__28207));
    LocalMux I__4638 (
            .O(N__28213),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv12 I__4637 (
            .O(N__28210),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__4636 (
            .O(N__28207),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__4635 (
            .O(N__28200),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__4634 (
            .O(N__28197),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__4633 (
            .O(N__28194),
            .I(N__28190));
    InMux I__4632 (
            .O(N__28193),
            .I(N__28186));
    LocalMux I__4631 (
            .O(N__28190),
            .I(N__28183));
    InMux I__4630 (
            .O(N__28189),
            .I(N__28180));
    LocalMux I__4629 (
            .O(N__28186),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv12 I__4628 (
            .O(N__28183),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__4627 (
            .O(N__28180),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__4626 (
            .O(N__28173),
            .I(N__28170));
    LocalMux I__4625 (
            .O(N__28170),
            .I(N__28167));
    Span4Mux_s2_v I__4624 (
            .O(N__28167),
            .I(N__28164));
    Odrv4 I__4623 (
            .O(N__28164),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    InMux I__4622 (
            .O(N__28161),
            .I(N__28156));
    InMux I__4621 (
            .O(N__28160),
            .I(N__28151));
    InMux I__4620 (
            .O(N__28159),
            .I(N__28151));
    LocalMux I__4619 (
            .O(N__28156),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__4618 (
            .O(N__28151),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    CascadeMux I__4617 (
            .O(N__28146),
            .I(N__28142));
    InMux I__4616 (
            .O(N__28145),
            .I(N__28138));
    InMux I__4615 (
            .O(N__28142),
            .I(N__28133));
    InMux I__4614 (
            .O(N__28141),
            .I(N__28133));
    LocalMux I__4613 (
            .O(N__28138),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__4612 (
            .O(N__28133),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    CascadeMux I__4611 (
            .O(N__28128),
            .I(N__28125));
    InMux I__4610 (
            .O(N__28125),
            .I(N__28122));
    LocalMux I__4609 (
            .O(N__28122),
            .I(N__28119));
    Span4Mux_h I__4608 (
            .O(N__28119),
            .I(N__28116));
    Odrv4 I__4607 (
            .O(N__28116),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    InMux I__4606 (
            .O(N__28113),
            .I(bfn_9_5_0_));
    InMux I__4605 (
            .O(N__28110),
            .I(N__28106));
    InMux I__4604 (
            .O(N__28109),
            .I(N__28103));
    LocalMux I__4603 (
            .O(N__28106),
            .I(N__28099));
    LocalMux I__4602 (
            .O(N__28103),
            .I(N__28096));
    InMux I__4601 (
            .O(N__28102),
            .I(N__28093));
    Span4Mux_v I__4600 (
            .O(N__28099),
            .I(N__28090));
    Span4Mux_h I__4599 (
            .O(N__28096),
            .I(N__28087));
    LocalMux I__4598 (
            .O(N__28093),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__4597 (
            .O(N__28090),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__4596 (
            .O(N__28087),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__4595 (
            .O(N__28080),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__4594 (
            .O(N__28077),
            .I(N__28072));
    InMux I__4593 (
            .O(N__28076),
            .I(N__28069));
    InMux I__4592 (
            .O(N__28075),
            .I(N__28066));
    LocalMux I__4591 (
            .O(N__28072),
            .I(N__28061));
    LocalMux I__4590 (
            .O(N__28069),
            .I(N__28061));
    LocalMux I__4589 (
            .O(N__28066),
            .I(N__28056));
    Span4Mux_v I__4588 (
            .O(N__28061),
            .I(N__28056));
    Odrv4 I__4587 (
            .O(N__28056),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__4586 (
            .O(N__28053),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__4585 (
            .O(N__28050),
            .I(N__28043));
    InMux I__4584 (
            .O(N__28049),
            .I(N__28043));
    InMux I__4583 (
            .O(N__28048),
            .I(N__28040));
    LocalMux I__4582 (
            .O(N__28043),
            .I(N__28037));
    LocalMux I__4581 (
            .O(N__28040),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__4580 (
            .O(N__28037),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__4579 (
            .O(N__28032),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    CascadeMux I__4578 (
            .O(N__28029),
            .I(N__28025));
    CascadeMux I__4577 (
            .O(N__28028),
            .I(N__28021));
    InMux I__4576 (
            .O(N__28025),
            .I(N__28016));
    InMux I__4575 (
            .O(N__28024),
            .I(N__28016));
    InMux I__4574 (
            .O(N__28021),
            .I(N__28013));
    LocalMux I__4573 (
            .O(N__28016),
            .I(N__28010));
    LocalMux I__4572 (
            .O(N__28013),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__4571 (
            .O(N__28010),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__4570 (
            .O(N__28005),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__4569 (
            .O(N__28002),
            .I(N__27997));
    InMux I__4568 (
            .O(N__28001),
            .I(N__27992));
    InMux I__4567 (
            .O(N__28000),
            .I(N__27992));
    LocalMux I__4566 (
            .O(N__27997),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    LocalMux I__4565 (
            .O(N__27992),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__4564 (
            .O(N__27987),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__4563 (
            .O(N__27984),
            .I(N__27979));
    InMux I__4562 (
            .O(N__27983),
            .I(N__27974));
    InMux I__4561 (
            .O(N__27982),
            .I(N__27974));
    LocalMux I__4560 (
            .O(N__27979),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    LocalMux I__4559 (
            .O(N__27974),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__4558 (
            .O(N__27969),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__4557 (
            .O(N__27966),
            .I(N__27961));
    InMux I__4556 (
            .O(N__27965),
            .I(N__27956));
    InMux I__4555 (
            .O(N__27964),
            .I(N__27956));
    LocalMux I__4554 (
            .O(N__27961),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    LocalMux I__4553 (
            .O(N__27956),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__4552 (
            .O(N__27951),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__4551 (
            .O(N__27948),
            .I(N__27943));
    InMux I__4550 (
            .O(N__27947),
            .I(N__27938));
    InMux I__4549 (
            .O(N__27946),
            .I(N__27938));
    LocalMux I__4548 (
            .O(N__27943),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    LocalMux I__4547 (
            .O(N__27938),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__4546 (
            .O(N__27933),
            .I(bfn_9_6_0_));
    InMux I__4545 (
            .O(N__27930),
            .I(N__27926));
    InMux I__4544 (
            .O(N__27929),
            .I(N__27923));
    LocalMux I__4543 (
            .O(N__27926),
            .I(N__27920));
    LocalMux I__4542 (
            .O(N__27923),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__4541 (
            .O(N__27920),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__4540 (
            .O(N__27915),
            .I(bfn_9_4_0_));
    InMux I__4539 (
            .O(N__27912),
            .I(N__27908));
    InMux I__4538 (
            .O(N__27911),
            .I(N__27905));
    LocalMux I__4537 (
            .O(N__27908),
            .I(N__27902));
    LocalMux I__4536 (
            .O(N__27905),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__4535 (
            .O(N__27902),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__4534 (
            .O(N__27897),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__4533 (
            .O(N__27894),
            .I(N__27890));
    InMux I__4532 (
            .O(N__27893),
            .I(N__27887));
    LocalMux I__4531 (
            .O(N__27890),
            .I(N__27884));
    LocalMux I__4530 (
            .O(N__27887),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__4529 (
            .O(N__27884),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__4528 (
            .O(N__27879),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__4527 (
            .O(N__27876),
            .I(N__27872));
    InMux I__4526 (
            .O(N__27875),
            .I(N__27869));
    LocalMux I__4525 (
            .O(N__27872),
            .I(N__27866));
    LocalMux I__4524 (
            .O(N__27869),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__4523 (
            .O(N__27866),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__4522 (
            .O(N__27861),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__4521 (
            .O(N__27858),
            .I(N__27855));
    LocalMux I__4520 (
            .O(N__27855),
            .I(N__27851));
    InMux I__4519 (
            .O(N__27854),
            .I(N__27848));
    Span4Mux_s1_v I__4518 (
            .O(N__27851),
            .I(N__27845));
    LocalMux I__4517 (
            .O(N__27848),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__4516 (
            .O(N__27845),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__4515 (
            .O(N__27840),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__4514 (
            .O(N__27837),
            .I(N__27834));
    LocalMux I__4513 (
            .O(N__27834),
            .I(N__27830));
    InMux I__4512 (
            .O(N__27833),
            .I(N__27827));
    Span4Mux_s1_v I__4511 (
            .O(N__27830),
            .I(N__27824));
    LocalMux I__4510 (
            .O(N__27827),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__4509 (
            .O(N__27824),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__4508 (
            .O(N__27819),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__4507 (
            .O(N__27816),
            .I(N__27812));
    InMux I__4506 (
            .O(N__27815),
            .I(N__27809));
    LocalMux I__4505 (
            .O(N__27812),
            .I(N__27806));
    LocalMux I__4504 (
            .O(N__27809),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__4503 (
            .O(N__27806),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__4502 (
            .O(N__27801),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__4501 (
            .O(N__27798),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__4500 (
            .O(N__27795),
            .I(N__27792));
    LocalMux I__4499 (
            .O(N__27792),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__4498 (
            .O(N__27789),
            .I(N__27785));
    CascadeMux I__4497 (
            .O(N__27788),
            .I(N__27782));
    InMux I__4496 (
            .O(N__27785),
            .I(N__27779));
    InMux I__4495 (
            .O(N__27782),
            .I(N__27775));
    LocalMux I__4494 (
            .O(N__27779),
            .I(N__27772));
    InMux I__4493 (
            .O(N__27778),
            .I(N__27769));
    LocalMux I__4492 (
            .O(N__27775),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__4491 (
            .O(N__27772),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__4490 (
            .O(N__27769),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__4489 (
            .O(N__27762),
            .I(N__27758));
    InMux I__4488 (
            .O(N__27761),
            .I(N__27755));
    LocalMux I__4487 (
            .O(N__27758),
            .I(N__27752));
    LocalMux I__4486 (
            .O(N__27755),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__4485 (
            .O(N__27752),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__4484 (
            .O(N__27747),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__4483 (
            .O(N__27744),
            .I(N__27740));
    InMux I__4482 (
            .O(N__27743),
            .I(N__27737));
    LocalMux I__4481 (
            .O(N__27740),
            .I(N__27734));
    LocalMux I__4480 (
            .O(N__27737),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__4479 (
            .O(N__27734),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__4478 (
            .O(N__27729),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__4477 (
            .O(N__27726),
            .I(N__27722));
    InMux I__4476 (
            .O(N__27725),
            .I(N__27719));
    LocalMux I__4475 (
            .O(N__27722),
            .I(N__27716));
    LocalMux I__4474 (
            .O(N__27719),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__4473 (
            .O(N__27716),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__4472 (
            .O(N__27711),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__4471 (
            .O(N__27708),
            .I(N__27704));
    InMux I__4470 (
            .O(N__27707),
            .I(N__27701));
    LocalMux I__4469 (
            .O(N__27704),
            .I(N__27698));
    LocalMux I__4468 (
            .O(N__27701),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__4467 (
            .O(N__27698),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__4466 (
            .O(N__27693),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__4465 (
            .O(N__27690),
            .I(N__27686));
    InMux I__4464 (
            .O(N__27689),
            .I(N__27683));
    LocalMux I__4463 (
            .O(N__27686),
            .I(N__27680));
    LocalMux I__4462 (
            .O(N__27683),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__4461 (
            .O(N__27680),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__4460 (
            .O(N__27675),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__4459 (
            .O(N__27672),
            .I(N__27669));
    LocalMux I__4458 (
            .O(N__27669),
            .I(N__27665));
    InMux I__4457 (
            .O(N__27668),
            .I(N__27662));
    Span4Mux_s1_v I__4456 (
            .O(N__27665),
            .I(N__27659));
    LocalMux I__4455 (
            .O(N__27662),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__4454 (
            .O(N__27659),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__4453 (
            .O(N__27654),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__4452 (
            .O(N__27651),
            .I(N__27647));
    InMux I__4451 (
            .O(N__27650),
            .I(N__27644));
    LocalMux I__4450 (
            .O(N__27647),
            .I(N__27641));
    LocalMux I__4449 (
            .O(N__27644),
            .I(N__27636));
    Span4Mux_s2_v I__4448 (
            .O(N__27641),
            .I(N__27636));
    Odrv4 I__4447 (
            .O(N__27636),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__4446 (
            .O(N__27633),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__4445 (
            .O(N__27630),
            .I(N__27626));
    InMux I__4444 (
            .O(N__27629),
            .I(N__27622));
    LocalMux I__4443 (
            .O(N__27626),
            .I(N__27619));
    InMux I__4442 (
            .O(N__27625),
            .I(N__27616));
    LocalMux I__4441 (
            .O(N__27622),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__4440 (
            .O(N__27619),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__4439 (
            .O(N__27616),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__4438 (
            .O(N__27609),
            .I(N__27605));
    InMux I__4437 (
            .O(N__27608),
            .I(N__27601));
    LocalMux I__4436 (
            .O(N__27605),
            .I(N__27598));
    InMux I__4435 (
            .O(N__27604),
            .I(N__27595));
    LocalMux I__4434 (
            .O(N__27601),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__4433 (
            .O(N__27598),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__4432 (
            .O(N__27595),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__4431 (
            .O(N__27588),
            .I(N__27583));
    InMux I__4430 (
            .O(N__27587),
            .I(N__27580));
    InMux I__4429 (
            .O(N__27586),
            .I(N__27577));
    LocalMux I__4428 (
            .O(N__27583),
            .I(N__27574));
    LocalMux I__4427 (
            .O(N__27580),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__4426 (
            .O(N__27577),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__4425 (
            .O(N__27574),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__4424 (
            .O(N__27567),
            .I(N__27564));
    LocalMux I__4423 (
            .O(N__27564),
            .I(N__27559));
    InMux I__4422 (
            .O(N__27563),
            .I(N__27556));
    InMux I__4421 (
            .O(N__27562),
            .I(N__27553));
    Span4Mux_v I__4420 (
            .O(N__27559),
            .I(N__27550));
    LocalMux I__4419 (
            .O(N__27556),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__4418 (
            .O(N__27553),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__4417 (
            .O(N__27550),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__4416 (
            .O(N__27543),
            .I(N__27539));
    InMux I__4415 (
            .O(N__27542),
            .I(N__27535));
    LocalMux I__4414 (
            .O(N__27539),
            .I(N__27532));
    InMux I__4413 (
            .O(N__27538),
            .I(N__27529));
    LocalMux I__4412 (
            .O(N__27535),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__4411 (
            .O(N__27532),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__4410 (
            .O(N__27529),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__4409 (
            .O(N__27522),
            .I(N__27517));
    InMux I__4408 (
            .O(N__27521),
            .I(N__27514));
    InMux I__4407 (
            .O(N__27520),
            .I(N__27511));
    LocalMux I__4406 (
            .O(N__27517),
            .I(N__27508));
    LocalMux I__4405 (
            .O(N__27514),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__4404 (
            .O(N__27511),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__4403 (
            .O(N__27508),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__4402 (
            .O(N__27501),
            .I(N__27496));
    InMux I__4401 (
            .O(N__27500),
            .I(N__27493));
    InMux I__4400 (
            .O(N__27499),
            .I(N__27490));
    LocalMux I__4399 (
            .O(N__27496),
            .I(N__27487));
    LocalMux I__4398 (
            .O(N__27493),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__4397 (
            .O(N__27490),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__4396 (
            .O(N__27487),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    CascadeMux I__4395 (
            .O(N__27480),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__4394 (
            .O(N__27477),
            .I(N__27472));
    InMux I__4393 (
            .O(N__27476),
            .I(N__27469));
    InMux I__4392 (
            .O(N__27475),
            .I(N__27466));
    LocalMux I__4391 (
            .O(N__27472),
            .I(N__27463));
    LocalMux I__4390 (
            .O(N__27469),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__4389 (
            .O(N__27466),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__4388 (
            .O(N__27463),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__4387 (
            .O(N__27456),
            .I(N__27453));
    LocalMux I__4386 (
            .O(N__27453),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__4385 (
            .O(N__27450),
            .I(N__27445));
    InMux I__4384 (
            .O(N__27449),
            .I(N__27442));
    InMux I__4383 (
            .O(N__27448),
            .I(N__27439));
    LocalMux I__4382 (
            .O(N__27445),
            .I(N__27436));
    LocalMux I__4381 (
            .O(N__27442),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__4380 (
            .O(N__27439),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__4379 (
            .O(N__27436),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    CascadeMux I__4378 (
            .O(N__27429),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__4377 (
            .O(N__27426),
            .I(N__27421));
    InMux I__4376 (
            .O(N__27425),
            .I(N__27418));
    InMux I__4375 (
            .O(N__27424),
            .I(N__27415));
    LocalMux I__4374 (
            .O(N__27421),
            .I(N__27412));
    LocalMux I__4373 (
            .O(N__27418),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__4372 (
            .O(N__27415),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__4371 (
            .O(N__27412),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__4370 (
            .O(N__27405),
            .I(N__27393));
    InMux I__4369 (
            .O(N__27404),
            .I(N__27393));
    InMux I__4368 (
            .O(N__27403),
            .I(N__27393));
    InMux I__4367 (
            .O(N__27402),
            .I(N__27393));
    LocalMux I__4366 (
            .O(N__27393),
            .I(N__27384));
    InMux I__4365 (
            .O(N__27392),
            .I(N__27379));
    InMux I__4364 (
            .O(N__27391),
            .I(N__27379));
    InMux I__4363 (
            .O(N__27390),
            .I(N__27370));
    InMux I__4362 (
            .O(N__27389),
            .I(N__27370));
    InMux I__4361 (
            .O(N__27388),
            .I(N__27370));
    InMux I__4360 (
            .O(N__27387),
            .I(N__27370));
    Odrv4 I__4359 (
            .O(N__27384),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__4358 (
            .O(N__27379),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__4357 (
            .O(N__27370),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__4356 (
            .O(N__27363),
            .I(N__27360));
    LocalMux I__4355 (
            .O(N__27360),
            .I(N__27357));
    Glb2LocalMux I__4354 (
            .O(N__27357),
            .I(N__27354));
    GlobalMux I__4353 (
            .O(N__27354),
            .I(clk_12mhz));
    IoInMux I__4352 (
            .O(N__27351),
            .I(N__27348));
    LocalMux I__4351 (
            .O(N__27348),
            .I(N__27345));
    IoSpan4Mux I__4350 (
            .O(N__27345),
            .I(N__27342));
    Odrv4 I__4349 (
            .O(N__27342),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__4348 (
            .O(N__27339),
            .I(N__27336));
    LocalMux I__4347 (
            .O(N__27336),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__4346 (
            .O(N__27333),
            .I(N__27330));
    LocalMux I__4345 (
            .O(N__27330),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__4344 (
            .O(N__27327),
            .I(N__27324));
    InMux I__4343 (
            .O(N__27324),
            .I(N__27321));
    LocalMux I__4342 (
            .O(N__27321),
            .I(\pwm_generator_inst.threshold_3 ));
    InMux I__4341 (
            .O(N__27318),
            .I(N__27315));
    LocalMux I__4340 (
            .O(N__27315),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__4339 (
            .O(N__27312),
            .I(N__27309));
    InMux I__4338 (
            .O(N__27309),
            .I(N__27306));
    LocalMux I__4337 (
            .O(N__27306),
            .I(N__27303));
    Sp12to4 I__4336 (
            .O(N__27303),
            .I(N__27300));
    Odrv12 I__4335 (
            .O(N__27300),
            .I(\pwm_generator_inst.threshold_4 ));
    InMux I__4334 (
            .O(N__27297),
            .I(N__27294));
    LocalMux I__4333 (
            .O(N__27294),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__4332 (
            .O(N__27291),
            .I(N__27288));
    InMux I__4331 (
            .O(N__27288),
            .I(N__27285));
    LocalMux I__4330 (
            .O(N__27285),
            .I(N__27282));
    Span4Mux_h I__4329 (
            .O(N__27282),
            .I(N__27279));
    Odrv4 I__4328 (
            .O(N__27279),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__4327 (
            .O(N__27276),
            .I(N__27273));
    LocalMux I__4326 (
            .O(N__27273),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__4325 (
            .O(N__27270),
            .I(N__27267));
    InMux I__4324 (
            .O(N__27267),
            .I(N__27264));
    LocalMux I__4323 (
            .O(N__27264),
            .I(\pwm_generator_inst.threshold_6 ));
    InMux I__4322 (
            .O(N__27261),
            .I(N__27258));
    LocalMux I__4321 (
            .O(N__27258),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__4320 (
            .O(N__27255),
            .I(N__27252));
    InMux I__4319 (
            .O(N__27252),
            .I(N__27249));
    LocalMux I__4318 (
            .O(N__27249),
            .I(\pwm_generator_inst.threshold_7 ));
    InMux I__4317 (
            .O(N__27246),
            .I(N__27243));
    LocalMux I__4316 (
            .O(N__27243),
            .I(N__27240));
    Odrv4 I__4315 (
            .O(N__27240),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__4314 (
            .O(N__27237),
            .I(N__27234));
    InMux I__4313 (
            .O(N__27234),
            .I(N__27231));
    LocalMux I__4312 (
            .O(N__27231),
            .I(\pwm_generator_inst.threshold_8 ));
    InMux I__4311 (
            .O(N__27228),
            .I(N__27225));
    LocalMux I__4310 (
            .O(N__27225),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__4309 (
            .O(N__27222),
            .I(N__27219));
    InMux I__4308 (
            .O(N__27219),
            .I(N__27216));
    LocalMux I__4307 (
            .O(N__27216),
            .I(N__27213));
    Odrv12 I__4306 (
            .O(N__27213),
            .I(\pwm_generator_inst.threshold_9 ));
    InMux I__4305 (
            .O(N__27210),
            .I(N__27207));
    LocalMux I__4304 (
            .O(N__27207),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__4303 (
            .O(N__27204),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__4302 (
            .O(N__27201),
            .I(N__27198));
    LocalMux I__4301 (
            .O(N__27198),
            .I(N__27195));
    IoSpan4Mux I__4300 (
            .O(N__27195),
            .I(N__27192));
    Span4Mux_s0_v I__4299 (
            .O(N__27192),
            .I(N__27189));
    Sp12to4 I__4298 (
            .O(N__27189),
            .I(N__27186));
    Span12Mux_v I__4297 (
            .O(N__27186),
            .I(N__27183));
    Span12Mux_h I__4296 (
            .O(N__27183),
            .I(N__27180));
    Odrv12 I__4295 (
            .O(N__27180),
            .I(pwm_output_c));
    CascadeMux I__4294 (
            .O(N__27177),
            .I(N__27174));
    InMux I__4293 (
            .O(N__27174),
            .I(N__27169));
    InMux I__4292 (
            .O(N__27173),
            .I(N__27166));
    InMux I__4291 (
            .O(N__27172),
            .I(N__27163));
    LocalMux I__4290 (
            .O(N__27169),
            .I(N__27158));
    LocalMux I__4289 (
            .O(N__27166),
            .I(N__27158));
    LocalMux I__4288 (
            .O(N__27163),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__4287 (
            .O(N__27158),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__4286 (
            .O(N__27153),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__4285 (
            .O(N__27150),
            .I(N__27146));
    InMux I__4284 (
            .O(N__27149),
            .I(N__27143));
    LocalMux I__4283 (
            .O(N__27146),
            .I(N__27140));
    LocalMux I__4282 (
            .O(N__27143),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv4 I__4281 (
            .O(N__27140),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__4280 (
            .O(N__27135),
            .I(N__27132));
    InMux I__4279 (
            .O(N__27132),
            .I(N__27127));
    InMux I__4278 (
            .O(N__27131),
            .I(N__27124));
    InMux I__4277 (
            .O(N__27130),
            .I(N__27121));
    LocalMux I__4276 (
            .O(N__27127),
            .I(N__27116));
    LocalMux I__4275 (
            .O(N__27124),
            .I(N__27116));
    LocalMux I__4274 (
            .O(N__27121),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__4273 (
            .O(N__27116),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__4272 (
            .O(N__27111),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__4271 (
            .O(N__27108),
            .I(N__27104));
    InMux I__4270 (
            .O(N__27107),
            .I(N__27101));
    LocalMux I__4269 (
            .O(N__27104),
            .I(N__27098));
    LocalMux I__4268 (
            .O(N__27101),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__4267 (
            .O(N__27098),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__4266 (
            .O(N__27093),
            .I(N__27090));
    InMux I__4265 (
            .O(N__27090),
            .I(N__27085));
    InMux I__4264 (
            .O(N__27089),
            .I(N__27082));
    InMux I__4263 (
            .O(N__27088),
            .I(N__27079));
    LocalMux I__4262 (
            .O(N__27085),
            .I(N__27074));
    LocalMux I__4261 (
            .O(N__27082),
            .I(N__27074));
    LocalMux I__4260 (
            .O(N__27079),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__4259 (
            .O(N__27074),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__4258 (
            .O(N__27069),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__4257 (
            .O(N__27066),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__4256 (
            .O(N__27063),
            .I(N__27056));
    CEMux I__4255 (
            .O(N__27062),
            .I(N__27053));
    CEMux I__4254 (
            .O(N__27061),
            .I(N__27050));
    CEMux I__4253 (
            .O(N__27060),
            .I(N__27047));
    CEMux I__4252 (
            .O(N__27059),
            .I(N__27044));
    LocalMux I__4251 (
            .O(N__27056),
            .I(N__27041));
    LocalMux I__4250 (
            .O(N__27053),
            .I(N__27038));
    LocalMux I__4249 (
            .O(N__27050),
            .I(N__27035));
    LocalMux I__4248 (
            .O(N__27047),
            .I(N__27032));
    LocalMux I__4247 (
            .O(N__27044),
            .I(N__27029));
    Span4Mux_v I__4246 (
            .O(N__27041),
            .I(N__27026));
    Span4Mux_v I__4245 (
            .O(N__27038),
            .I(N__27023));
    Span4Mux_v I__4244 (
            .O(N__27035),
            .I(N__27020));
    Span4Mux_v I__4243 (
            .O(N__27032),
            .I(N__27015));
    Span4Mux_v I__4242 (
            .O(N__27029),
            .I(N__27015));
    Odrv4 I__4241 (
            .O(N__27026),
            .I(\delay_measurement_inst.delay_tr_timer.N_165_i ));
    Odrv4 I__4240 (
            .O(N__27023),
            .I(\delay_measurement_inst.delay_tr_timer.N_165_i ));
    Odrv4 I__4239 (
            .O(N__27020),
            .I(\delay_measurement_inst.delay_tr_timer.N_165_i ));
    Odrv4 I__4238 (
            .O(N__27015),
            .I(\delay_measurement_inst.delay_tr_timer.N_165_i ));
    InMux I__4237 (
            .O(N__27006),
            .I(N__26991));
    InMux I__4236 (
            .O(N__27005),
            .I(N__26991));
    InMux I__4235 (
            .O(N__27004),
            .I(N__26991));
    InMux I__4234 (
            .O(N__27003),
            .I(N__26991));
    InMux I__4233 (
            .O(N__27002),
            .I(N__26991));
    LocalMux I__4232 (
            .O(N__26991),
            .I(N__26985));
    InMux I__4231 (
            .O(N__26990),
            .I(N__26980));
    InMux I__4230 (
            .O(N__26989),
            .I(N__26977));
    InMux I__4229 (
            .O(N__26988),
            .I(N__26974));
    Span4Mux_h I__4228 (
            .O(N__26985),
            .I(N__26971));
    InMux I__4227 (
            .O(N__26984),
            .I(N__26966));
    InMux I__4226 (
            .O(N__26983),
            .I(N__26966));
    LocalMux I__4225 (
            .O(N__26980),
            .I(N__26963));
    LocalMux I__4224 (
            .O(N__26977),
            .I(N__26960));
    LocalMux I__4223 (
            .O(N__26974),
            .I(N__26957));
    Span4Mux_v I__4222 (
            .O(N__26971),
            .I(N__26952));
    LocalMux I__4221 (
            .O(N__26966),
            .I(N__26952));
    Span12Mux_h I__4220 (
            .O(N__26963),
            .I(N__26949));
    Span4Mux_v I__4219 (
            .O(N__26960),
            .I(N__26944));
    Span4Mux_h I__4218 (
            .O(N__26957),
            .I(N__26944));
    Span4Mux_h I__4217 (
            .O(N__26952),
            .I(N__26941));
    Odrv12 I__4216 (
            .O(N__26949),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__4215 (
            .O(N__26944),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__4214 (
            .O(N__26941),
            .I(\pwm_generator_inst.N_16 ));
    InMux I__4213 (
            .O(N__26934),
            .I(N__26931));
    LocalMux I__4212 (
            .O(N__26931),
            .I(N__26928));
    Span4Mux_v I__4211 (
            .O(N__26928),
            .I(N__26925));
    Span4Mux_h I__4210 (
            .O(N__26925),
            .I(N__26922));
    Odrv4 I__4209 (
            .O(N__26922),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ));
    InMux I__4208 (
            .O(N__26919),
            .I(N__26908));
    InMux I__4207 (
            .O(N__26918),
            .I(N__26903));
    InMux I__4206 (
            .O(N__26917),
            .I(N__26903));
    InMux I__4205 (
            .O(N__26916),
            .I(N__26900));
    InMux I__4204 (
            .O(N__26915),
            .I(N__26889));
    InMux I__4203 (
            .O(N__26914),
            .I(N__26889));
    InMux I__4202 (
            .O(N__26913),
            .I(N__26889));
    InMux I__4201 (
            .O(N__26912),
            .I(N__26889));
    InMux I__4200 (
            .O(N__26911),
            .I(N__26889));
    LocalMux I__4199 (
            .O(N__26908),
            .I(N__26884));
    LocalMux I__4198 (
            .O(N__26903),
            .I(N__26884));
    LocalMux I__4197 (
            .O(N__26900),
            .I(N__26879));
    LocalMux I__4196 (
            .O(N__26889),
            .I(N__26879));
    Span4Mux_v I__4195 (
            .O(N__26884),
            .I(N__26875));
    Span4Mux_v I__4194 (
            .O(N__26879),
            .I(N__26872));
    InMux I__4193 (
            .O(N__26878),
            .I(N__26869));
    Sp12to4 I__4192 (
            .O(N__26875),
            .I(N__26862));
    Sp12to4 I__4191 (
            .O(N__26872),
            .I(N__26862));
    LocalMux I__4190 (
            .O(N__26869),
            .I(N__26862));
    Odrv12 I__4189 (
            .O(N__26862),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__4188 (
            .O(N__26859),
            .I(N__26856));
    InMux I__4187 (
            .O(N__26856),
            .I(N__26853));
    LocalMux I__4186 (
            .O(N__26853),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__4185 (
            .O(N__26850),
            .I(N__26847));
    LocalMux I__4184 (
            .O(N__26847),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__4183 (
            .O(N__26844),
            .I(N__26841));
    InMux I__4182 (
            .O(N__26841),
            .I(N__26838));
    LocalMux I__4181 (
            .O(N__26838),
            .I(N__26835));
    Odrv4 I__4180 (
            .O(N__26835),
            .I(\pwm_generator_inst.threshold_1 ));
    InMux I__4179 (
            .O(N__26832),
            .I(N__26829));
    LocalMux I__4178 (
            .O(N__26829),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__4177 (
            .O(N__26826),
            .I(N__26823));
    InMux I__4176 (
            .O(N__26823),
            .I(N__26820));
    LocalMux I__4175 (
            .O(N__26820),
            .I(N__26817));
    Odrv12 I__4174 (
            .O(N__26817),
            .I(\pwm_generator_inst.threshold_2 ));
    InMux I__4173 (
            .O(N__26814),
            .I(N__26811));
    LocalMux I__4172 (
            .O(N__26811),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__4171 (
            .O(N__26808),
            .I(N__26805));
    InMux I__4170 (
            .O(N__26805),
            .I(N__26800));
    InMux I__4169 (
            .O(N__26804),
            .I(N__26797));
    InMux I__4168 (
            .O(N__26803),
            .I(N__26794));
    LocalMux I__4167 (
            .O(N__26800),
            .I(N__26789));
    LocalMux I__4166 (
            .O(N__26797),
            .I(N__26789));
    LocalMux I__4165 (
            .O(N__26794),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__4164 (
            .O(N__26789),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__4163 (
            .O(N__26784),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__4162 (
            .O(N__26781),
            .I(N__26774));
    InMux I__4161 (
            .O(N__26780),
            .I(N__26774));
    InMux I__4160 (
            .O(N__26779),
            .I(N__26771));
    LocalMux I__4159 (
            .O(N__26774),
            .I(N__26768));
    LocalMux I__4158 (
            .O(N__26771),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__4157 (
            .O(N__26768),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__4156 (
            .O(N__26763),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__4155 (
            .O(N__26760),
            .I(N__26753));
    InMux I__4154 (
            .O(N__26759),
            .I(N__26753));
    InMux I__4153 (
            .O(N__26758),
            .I(N__26750));
    LocalMux I__4152 (
            .O(N__26753),
            .I(N__26747));
    LocalMux I__4151 (
            .O(N__26750),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__4150 (
            .O(N__26747),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__4149 (
            .O(N__26742),
            .I(N__26737));
    InMux I__4148 (
            .O(N__26741),
            .I(N__26732));
    InMux I__4147 (
            .O(N__26740),
            .I(N__26732));
    LocalMux I__4146 (
            .O(N__26737),
            .I(N__26728));
    LocalMux I__4145 (
            .O(N__26732),
            .I(N__26725));
    InMux I__4144 (
            .O(N__26731),
            .I(N__26722));
    Sp12to4 I__4143 (
            .O(N__26728),
            .I(N__26715));
    Span12Mux_s3_v I__4142 (
            .O(N__26725),
            .I(N__26715));
    LocalMux I__4141 (
            .O(N__26722),
            .I(N__26715));
    Odrv12 I__4140 (
            .O(N__26715),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__4139 (
            .O(N__26712),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__4138 (
            .O(N__26709),
            .I(N__26705));
    InMux I__4137 (
            .O(N__26708),
            .I(N__26702));
    InMux I__4136 (
            .O(N__26705),
            .I(N__26699));
    LocalMux I__4135 (
            .O(N__26702),
            .I(N__26693));
    LocalMux I__4134 (
            .O(N__26699),
            .I(N__26693));
    InMux I__4133 (
            .O(N__26698),
            .I(N__26690));
    Span4Mux_h I__4132 (
            .O(N__26693),
            .I(N__26687));
    LocalMux I__4131 (
            .O(N__26690),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__4130 (
            .O(N__26687),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    CascadeMux I__4129 (
            .O(N__26682),
            .I(N__26678));
    InMux I__4128 (
            .O(N__26681),
            .I(N__26673));
    InMux I__4127 (
            .O(N__26678),
            .I(N__26670));
    InMux I__4126 (
            .O(N__26677),
            .I(N__26667));
    InMux I__4125 (
            .O(N__26676),
            .I(N__26664));
    LocalMux I__4124 (
            .O(N__26673),
            .I(N__26661));
    LocalMux I__4123 (
            .O(N__26670),
            .I(N__26654));
    LocalMux I__4122 (
            .O(N__26667),
            .I(N__26654));
    LocalMux I__4121 (
            .O(N__26664),
            .I(N__26654));
    Span4Mux_h I__4120 (
            .O(N__26661),
            .I(N__26649));
    Span4Mux_v I__4119 (
            .O(N__26654),
            .I(N__26649));
    Odrv4 I__4118 (
            .O(N__26649),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__4117 (
            .O(N__26646),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__4116 (
            .O(N__26643),
            .I(N__26639));
    CascadeMux I__4115 (
            .O(N__26642),
            .I(N__26636));
    InMux I__4114 (
            .O(N__26639),
            .I(N__26631));
    InMux I__4113 (
            .O(N__26636),
            .I(N__26631));
    LocalMux I__4112 (
            .O(N__26631),
            .I(N__26627));
    InMux I__4111 (
            .O(N__26630),
            .I(N__26624));
    Span4Mux_h I__4110 (
            .O(N__26627),
            .I(N__26621));
    LocalMux I__4109 (
            .O(N__26624),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv4 I__4108 (
            .O(N__26621),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__4107 (
            .O(N__26616),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__4106 (
            .O(N__26613),
            .I(N__26609));
    CascadeMux I__4105 (
            .O(N__26612),
            .I(N__26606));
    InMux I__4104 (
            .O(N__26609),
            .I(N__26600));
    InMux I__4103 (
            .O(N__26606),
            .I(N__26600));
    InMux I__4102 (
            .O(N__26605),
            .I(N__26597));
    LocalMux I__4101 (
            .O(N__26600),
            .I(N__26594));
    LocalMux I__4100 (
            .O(N__26597),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__4099 (
            .O(N__26594),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__4098 (
            .O(N__26589),
            .I(N__26584));
    InMux I__4097 (
            .O(N__26588),
            .I(N__26579));
    InMux I__4096 (
            .O(N__26587),
            .I(N__26579));
    LocalMux I__4095 (
            .O(N__26584),
            .I(N__26575));
    LocalMux I__4094 (
            .O(N__26579),
            .I(N__26572));
    InMux I__4093 (
            .O(N__26578),
            .I(N__26569));
    Sp12to4 I__4092 (
            .O(N__26575),
            .I(N__26562));
    Span12Mux_s6_v I__4091 (
            .O(N__26572),
            .I(N__26562));
    LocalMux I__4090 (
            .O(N__26569),
            .I(N__26562));
    Odrv12 I__4089 (
            .O(N__26562),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__4088 (
            .O(N__26559),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__4087 (
            .O(N__26556),
            .I(N__26553));
    InMux I__4086 (
            .O(N__26553),
            .I(N__26549));
    InMux I__4085 (
            .O(N__26552),
            .I(N__26546));
    LocalMux I__4084 (
            .O(N__26549),
            .I(N__26540));
    LocalMux I__4083 (
            .O(N__26546),
            .I(N__26540));
    InMux I__4082 (
            .O(N__26545),
            .I(N__26537));
    Span4Mux_h I__4081 (
            .O(N__26540),
            .I(N__26534));
    LocalMux I__4080 (
            .O(N__26537),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__4079 (
            .O(N__26534),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__4078 (
            .O(N__26529),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__4077 (
            .O(N__26526),
            .I(N__26523));
    InMux I__4076 (
            .O(N__26523),
            .I(N__26518));
    InMux I__4075 (
            .O(N__26522),
            .I(N__26515));
    InMux I__4074 (
            .O(N__26521),
            .I(N__26512));
    LocalMux I__4073 (
            .O(N__26518),
            .I(N__26507));
    LocalMux I__4072 (
            .O(N__26515),
            .I(N__26507));
    LocalMux I__4071 (
            .O(N__26512),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__4070 (
            .O(N__26507),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__4069 (
            .O(N__26502),
            .I(bfn_8_14_0_));
    CascadeMux I__4068 (
            .O(N__26499),
            .I(N__26496));
    InMux I__4067 (
            .O(N__26496),
            .I(N__26493));
    LocalMux I__4066 (
            .O(N__26493),
            .I(N__26488));
    InMux I__4065 (
            .O(N__26492),
            .I(N__26485));
    InMux I__4064 (
            .O(N__26491),
            .I(N__26482));
    Span4Mux_h I__4063 (
            .O(N__26488),
            .I(N__26479));
    LocalMux I__4062 (
            .O(N__26485),
            .I(N__26476));
    LocalMux I__4061 (
            .O(N__26482),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__4060 (
            .O(N__26479),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__4059 (
            .O(N__26476),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__4058 (
            .O(N__26469),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__4057 (
            .O(N__26466),
            .I(N__26463));
    InMux I__4056 (
            .O(N__26463),
            .I(N__26458));
    InMux I__4055 (
            .O(N__26462),
            .I(N__26455));
    InMux I__4054 (
            .O(N__26461),
            .I(N__26452));
    LocalMux I__4053 (
            .O(N__26458),
            .I(N__26447));
    LocalMux I__4052 (
            .O(N__26455),
            .I(N__26447));
    LocalMux I__4051 (
            .O(N__26452),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__4050 (
            .O(N__26447),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__4049 (
            .O(N__26442),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__4048 (
            .O(N__26439),
            .I(N__26433));
    InMux I__4047 (
            .O(N__26438),
            .I(N__26433));
    LocalMux I__4046 (
            .O(N__26433),
            .I(N__26429));
    InMux I__4045 (
            .O(N__26432),
            .I(N__26426));
    Span4Mux_v I__4044 (
            .O(N__26429),
            .I(N__26423));
    LocalMux I__4043 (
            .O(N__26426),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__4042 (
            .O(N__26423),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__4041 (
            .O(N__26418),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__4040 (
            .O(N__26415),
            .I(N__26408));
    InMux I__4039 (
            .O(N__26414),
            .I(N__26408));
    InMux I__4038 (
            .O(N__26413),
            .I(N__26405));
    LocalMux I__4037 (
            .O(N__26408),
            .I(N__26402));
    LocalMux I__4036 (
            .O(N__26405),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__4035 (
            .O(N__26402),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__4034 (
            .O(N__26397),
            .I(N__26393));
    InMux I__4033 (
            .O(N__26396),
            .I(N__26390));
    LocalMux I__4032 (
            .O(N__26393),
            .I(N__26386));
    LocalMux I__4031 (
            .O(N__26390),
            .I(N__26383));
    InMux I__4030 (
            .O(N__26389),
            .I(N__26380));
    Span4Mux_h I__4029 (
            .O(N__26386),
            .I(N__26376));
    Span4Mux_s3_v I__4028 (
            .O(N__26383),
            .I(N__26371));
    LocalMux I__4027 (
            .O(N__26380),
            .I(N__26371));
    InMux I__4026 (
            .O(N__26379),
            .I(N__26368));
    Span4Mux_v I__4025 (
            .O(N__26376),
            .I(N__26365));
    Span4Mux_v I__4024 (
            .O(N__26371),
            .I(N__26360));
    LocalMux I__4023 (
            .O(N__26368),
            .I(N__26360));
    Odrv4 I__4022 (
            .O(N__26365),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv4 I__4021 (
            .O(N__26360),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__4020 (
            .O(N__26355),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__4019 (
            .O(N__26352),
            .I(N__26348));
    CascadeMux I__4018 (
            .O(N__26351),
            .I(N__26345));
    InMux I__4017 (
            .O(N__26348),
            .I(N__26339));
    InMux I__4016 (
            .O(N__26345),
            .I(N__26339));
    InMux I__4015 (
            .O(N__26344),
            .I(N__26336));
    LocalMux I__4014 (
            .O(N__26339),
            .I(N__26333));
    LocalMux I__4013 (
            .O(N__26336),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__4012 (
            .O(N__26333),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__4011 (
            .O(N__26328),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__4010 (
            .O(N__26325),
            .I(N__26321));
    CascadeMux I__4009 (
            .O(N__26324),
            .I(N__26318));
    InMux I__4008 (
            .O(N__26321),
            .I(N__26313));
    InMux I__4007 (
            .O(N__26318),
            .I(N__26313));
    LocalMux I__4006 (
            .O(N__26313),
            .I(N__26309));
    InMux I__4005 (
            .O(N__26312),
            .I(N__26306));
    Span4Mux_h I__4004 (
            .O(N__26309),
            .I(N__26303));
    LocalMux I__4003 (
            .O(N__26306),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__4002 (
            .O(N__26303),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__4001 (
            .O(N__26298),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__4000 (
            .O(N__26295),
            .I(N__26292));
    InMux I__3999 (
            .O(N__26292),
            .I(N__26287));
    InMux I__3998 (
            .O(N__26291),
            .I(N__26284));
    InMux I__3997 (
            .O(N__26290),
            .I(N__26281));
    LocalMux I__3996 (
            .O(N__26287),
            .I(N__26276));
    LocalMux I__3995 (
            .O(N__26284),
            .I(N__26276));
    LocalMux I__3994 (
            .O(N__26281),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__3993 (
            .O(N__26276),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__3992 (
            .O(N__26271),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__3991 (
            .O(N__26268),
            .I(N__26265));
    InMux I__3990 (
            .O(N__26265),
            .I(N__26260));
    InMux I__3989 (
            .O(N__26264),
            .I(N__26257));
    InMux I__3988 (
            .O(N__26263),
            .I(N__26254));
    LocalMux I__3987 (
            .O(N__26260),
            .I(N__26249));
    LocalMux I__3986 (
            .O(N__26257),
            .I(N__26249));
    LocalMux I__3985 (
            .O(N__26254),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__3984 (
            .O(N__26249),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__3983 (
            .O(N__26244),
            .I(bfn_8_13_0_));
    CascadeMux I__3982 (
            .O(N__26241),
            .I(N__26237));
    InMux I__3981 (
            .O(N__26240),
            .I(N__26234));
    InMux I__3980 (
            .O(N__26237),
            .I(N__26231));
    LocalMux I__3979 (
            .O(N__26234),
            .I(N__26225));
    LocalMux I__3978 (
            .O(N__26231),
            .I(N__26225));
    InMux I__3977 (
            .O(N__26230),
            .I(N__26222));
    Span4Mux_h I__3976 (
            .O(N__26225),
            .I(N__26219));
    LocalMux I__3975 (
            .O(N__26222),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__3974 (
            .O(N__26219),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__3973 (
            .O(N__26214),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__3972 (
            .O(N__26211),
            .I(N__26205));
    InMux I__3971 (
            .O(N__26210),
            .I(N__26205));
    LocalMux I__3970 (
            .O(N__26205),
            .I(N__26201));
    InMux I__3969 (
            .O(N__26204),
            .I(N__26198));
    Span4Mux_v I__3968 (
            .O(N__26201),
            .I(N__26195));
    LocalMux I__3967 (
            .O(N__26198),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__3966 (
            .O(N__26195),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__3965 (
            .O(N__26190),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__3964 (
            .O(N__26187),
            .I(N__26180));
    InMux I__3963 (
            .O(N__26186),
            .I(N__26180));
    InMux I__3962 (
            .O(N__26185),
            .I(N__26177));
    LocalMux I__3961 (
            .O(N__26180),
            .I(N__26174));
    LocalMux I__3960 (
            .O(N__26177),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__3959 (
            .O(N__26174),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__3958 (
            .O(N__26169),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__3957 (
            .O(N__26166),
            .I(N__26162));
    CascadeMux I__3956 (
            .O(N__26165),
            .I(N__26159));
    InMux I__3955 (
            .O(N__26162),
            .I(N__26153));
    InMux I__3954 (
            .O(N__26159),
            .I(N__26153));
    InMux I__3953 (
            .O(N__26158),
            .I(N__26150));
    LocalMux I__3952 (
            .O(N__26153),
            .I(N__26147));
    LocalMux I__3951 (
            .O(N__26150),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv4 I__3950 (
            .O(N__26147),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__3949 (
            .O(N__26142),
            .I(N__26137));
    InMux I__3948 (
            .O(N__26141),
            .I(N__26134));
    InMux I__3947 (
            .O(N__26140),
            .I(N__26131));
    LocalMux I__3946 (
            .O(N__26137),
            .I(N__26126));
    LocalMux I__3945 (
            .O(N__26134),
            .I(N__26126));
    LocalMux I__3944 (
            .O(N__26131),
            .I(N__26122));
    Sp12to4 I__3943 (
            .O(N__26126),
            .I(N__26119));
    InMux I__3942 (
            .O(N__26125),
            .I(N__26116));
    Odrv4 I__3941 (
            .O(N__26122),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv12 I__3940 (
            .O(N__26119),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    LocalMux I__3939 (
            .O(N__26116),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__3938 (
            .O(N__26109),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__3937 (
            .O(N__26106),
            .I(N__26102));
    CascadeMux I__3936 (
            .O(N__26105),
            .I(N__26099));
    InMux I__3935 (
            .O(N__26102),
            .I(N__26093));
    InMux I__3934 (
            .O(N__26099),
            .I(N__26093));
    InMux I__3933 (
            .O(N__26098),
            .I(N__26090));
    LocalMux I__3932 (
            .O(N__26093),
            .I(N__26087));
    LocalMux I__3931 (
            .O(N__26090),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__3930 (
            .O(N__26087),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__3929 (
            .O(N__26082),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__3928 (
            .O(N__26079),
            .I(N__26076));
    InMux I__3927 (
            .O(N__26076),
            .I(N__26071));
    InMux I__3926 (
            .O(N__26075),
            .I(N__26068));
    InMux I__3925 (
            .O(N__26074),
            .I(N__26065));
    LocalMux I__3924 (
            .O(N__26071),
            .I(N__26060));
    LocalMux I__3923 (
            .O(N__26068),
            .I(N__26060));
    LocalMux I__3922 (
            .O(N__26065),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__3921 (
            .O(N__26060),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__3920 (
            .O(N__26055),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__3919 (
            .O(N__26052),
            .I(N__26049));
    InMux I__3918 (
            .O(N__26049),
            .I(N__26045));
    InMux I__3917 (
            .O(N__26048),
            .I(N__26042));
    LocalMux I__3916 (
            .O(N__26045),
            .I(N__26036));
    LocalMux I__3915 (
            .O(N__26042),
            .I(N__26036));
    InMux I__3914 (
            .O(N__26041),
            .I(N__26033));
    Span4Mux_h I__3913 (
            .O(N__26036),
            .I(N__26030));
    LocalMux I__3912 (
            .O(N__26033),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__3911 (
            .O(N__26030),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__3910 (
            .O(N__26025),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__3909 (
            .O(N__26022),
            .I(N__26019));
    InMux I__3908 (
            .O(N__26019),
            .I(N__26014));
    InMux I__3907 (
            .O(N__26018),
            .I(N__26011));
    InMux I__3906 (
            .O(N__26017),
            .I(N__26008));
    LocalMux I__3905 (
            .O(N__26014),
            .I(N__26003));
    LocalMux I__3904 (
            .O(N__26011),
            .I(N__26003));
    LocalMux I__3903 (
            .O(N__26008),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__3902 (
            .O(N__26003),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__3901 (
            .O(N__25998),
            .I(N__25995));
    LocalMux I__3900 (
            .O(N__25995),
            .I(N__25990));
    InMux I__3899 (
            .O(N__25994),
            .I(N__25987));
    InMux I__3898 (
            .O(N__25993),
            .I(N__25983));
    Span4Mux_h I__3897 (
            .O(N__25990),
            .I(N__25980));
    LocalMux I__3896 (
            .O(N__25987),
            .I(N__25977));
    InMux I__3895 (
            .O(N__25986),
            .I(N__25974));
    LocalMux I__3894 (
            .O(N__25983),
            .I(N__25971));
    Span4Mux_v I__3893 (
            .O(N__25980),
            .I(N__25968));
    Sp12to4 I__3892 (
            .O(N__25977),
            .I(N__25963));
    LocalMux I__3891 (
            .O(N__25974),
            .I(N__25963));
    Odrv4 I__3890 (
            .O(N__25971),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    Odrv4 I__3889 (
            .O(N__25968),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    Odrv12 I__3888 (
            .O(N__25963),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__3887 (
            .O(N__25956),
            .I(bfn_8_12_0_));
    CascadeMux I__3886 (
            .O(N__25953),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    CascadeMux I__3885 (
            .O(N__25950),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ));
    InMux I__3884 (
            .O(N__25947),
            .I(N__25944));
    LocalMux I__3883 (
            .O(N__25944),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ));
    CascadeMux I__3882 (
            .O(N__25941),
            .I(N__25938));
    InMux I__3881 (
            .O(N__25938),
            .I(N__25935));
    LocalMux I__3880 (
            .O(N__25935),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ));
    CascadeMux I__3879 (
            .O(N__25932),
            .I(N__25928));
    InMux I__3878 (
            .O(N__25931),
            .I(N__25925));
    InMux I__3877 (
            .O(N__25928),
            .I(N__25922));
    LocalMux I__3876 (
            .O(N__25925),
            .I(N__25916));
    LocalMux I__3875 (
            .O(N__25922),
            .I(N__25916));
    InMux I__3874 (
            .O(N__25921),
            .I(N__25913));
    Span4Mux_h I__3873 (
            .O(N__25916),
            .I(N__25910));
    LocalMux I__3872 (
            .O(N__25913),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__3871 (
            .O(N__25910),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__3870 (
            .O(N__25905),
            .I(N__25902));
    LocalMux I__3869 (
            .O(N__25902),
            .I(N__25899));
    Span4Mux_s3_v I__3868 (
            .O(N__25899),
            .I(N__25896));
    Odrv4 I__3867 (
            .O(N__25896),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__3866 (
            .O(N__25893),
            .I(N__25890));
    InMux I__3865 (
            .O(N__25890),
            .I(N__25884));
    InMux I__3864 (
            .O(N__25889),
            .I(N__25884));
    LocalMux I__3863 (
            .O(N__25884),
            .I(N__25881));
    Span4Mux_h I__3862 (
            .O(N__25881),
            .I(N__25878));
    Odrv4 I__3861 (
            .O(N__25878),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    InMux I__3860 (
            .O(N__25875),
            .I(N__25870));
    InMux I__3859 (
            .O(N__25874),
            .I(N__25867));
    InMux I__3858 (
            .O(N__25873),
            .I(N__25864));
    LocalMux I__3857 (
            .O(N__25870),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__3856 (
            .O(N__25867),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__3855 (
            .O(N__25864),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__3854 (
            .O(N__25857),
            .I(N__25854));
    LocalMux I__3853 (
            .O(N__25854),
            .I(N__25851));
    Odrv4 I__3852 (
            .O(N__25851),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ));
    CascadeMux I__3851 (
            .O(N__25848),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ));
    InMux I__3850 (
            .O(N__25845),
            .I(N__25839));
    InMux I__3849 (
            .O(N__25844),
            .I(N__25839));
    LocalMux I__3848 (
            .O(N__25839),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    InMux I__3847 (
            .O(N__25836),
            .I(N__25833));
    LocalMux I__3846 (
            .O(N__25833),
            .I(N__25830));
    Odrv12 I__3845 (
            .O(N__25830),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__3844 (
            .O(N__25827),
            .I(N__25824));
    InMux I__3843 (
            .O(N__25824),
            .I(N__25821));
    LocalMux I__3842 (
            .O(N__25821),
            .I(N__25818));
    Odrv4 I__3841 (
            .O(N__25818),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    InMux I__3840 (
            .O(N__25815),
            .I(N__25812));
    LocalMux I__3839 (
            .O(N__25812),
            .I(N__25809));
    Odrv4 I__3838 (
            .O(N__25809),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    CascadeMux I__3837 (
            .O(N__25806),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_));
    CascadeMux I__3836 (
            .O(N__25803),
            .I(N__25800));
    InMux I__3835 (
            .O(N__25800),
            .I(N__25794));
    InMux I__3834 (
            .O(N__25799),
            .I(N__25794));
    LocalMux I__3833 (
            .O(N__25794),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    InMux I__3832 (
            .O(N__25791),
            .I(N__25785));
    InMux I__3831 (
            .O(N__25790),
            .I(N__25785));
    LocalMux I__3830 (
            .O(N__25785),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    InMux I__3829 (
            .O(N__25782),
            .I(N__25779));
    LocalMux I__3828 (
            .O(N__25779),
            .I(N__25776));
    Span4Mux_h I__3827 (
            .O(N__25776),
            .I(N__25772));
    InMux I__3826 (
            .O(N__25775),
            .I(N__25769));
    Odrv4 I__3825 (
            .O(N__25772),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    LocalMux I__3824 (
            .O(N__25769),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__3823 (
            .O(N__25764),
            .I(N__25760));
    CascadeMux I__3822 (
            .O(N__25763),
            .I(N__25757));
    InMux I__3821 (
            .O(N__25760),
            .I(N__25754));
    InMux I__3820 (
            .O(N__25757),
            .I(N__25751));
    LocalMux I__3819 (
            .O(N__25754),
            .I(N__25748));
    LocalMux I__3818 (
            .O(N__25751),
            .I(N__25745));
    Span4Mux_v I__3817 (
            .O(N__25748),
            .I(N__25742));
    Span4Mux_v I__3816 (
            .O(N__25745),
            .I(N__25739));
    Odrv4 I__3815 (
            .O(N__25742),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    Odrv4 I__3814 (
            .O(N__25739),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    InMux I__3813 (
            .O(N__25734),
            .I(N__25731));
    LocalMux I__3812 (
            .O(N__25731),
            .I(N__25728));
    Span4Mux_s3_v I__3811 (
            .O(N__25728),
            .I(N__25725));
    Odrv4 I__3810 (
            .O(N__25725),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ));
    InMux I__3809 (
            .O(N__25722),
            .I(N__25719));
    LocalMux I__3808 (
            .O(N__25719),
            .I(N__25716));
    Odrv12 I__3807 (
            .O(N__25716),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    InMux I__3806 (
            .O(N__25713),
            .I(N__25710));
    LocalMux I__3805 (
            .O(N__25710),
            .I(N__25707));
    Span4Mux_v I__3804 (
            .O(N__25707),
            .I(N__25703));
    InMux I__3803 (
            .O(N__25706),
            .I(N__25700));
    Odrv4 I__3802 (
            .O(N__25703),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__3801 (
            .O(N__25700),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    CascadeMux I__3800 (
            .O(N__25695),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_));
    InMux I__3799 (
            .O(N__25692),
            .I(N__25686));
    InMux I__3798 (
            .O(N__25691),
            .I(N__25686));
    LocalMux I__3797 (
            .O(N__25686),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    CascadeMux I__3796 (
            .O(N__25683),
            .I(N__25679));
    CascadeMux I__3795 (
            .O(N__25682),
            .I(N__25676));
    InMux I__3794 (
            .O(N__25679),
            .I(N__25671));
    InMux I__3793 (
            .O(N__25676),
            .I(N__25671));
    LocalMux I__3792 (
            .O(N__25671),
            .I(N__25668));
    Span4Mux_h I__3791 (
            .O(N__25668),
            .I(N__25665));
    Odrv4 I__3790 (
            .O(N__25665),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    InMux I__3789 (
            .O(N__25662),
            .I(N__25659));
    LocalMux I__3788 (
            .O(N__25659),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    InMux I__3787 (
            .O(N__25656),
            .I(N__25653));
    LocalMux I__3786 (
            .O(N__25653),
            .I(N__25650));
    Odrv12 I__3785 (
            .O(N__25650),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__3784 (
            .O(N__25647),
            .I(N__25644));
    InMux I__3783 (
            .O(N__25644),
            .I(N__25641));
    LocalMux I__3782 (
            .O(N__25641),
            .I(N__25638));
    Odrv4 I__3781 (
            .O(N__25638),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    InMux I__3780 (
            .O(N__25635),
            .I(N__25632));
    LocalMux I__3779 (
            .O(N__25632),
            .I(N__25629));
    Span4Mux_v I__3778 (
            .O(N__25629),
            .I(N__25625));
    InMux I__3777 (
            .O(N__25628),
            .I(N__25622));
    Odrv4 I__3776 (
            .O(N__25625),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    LocalMux I__3775 (
            .O(N__25622),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    CascadeMux I__3774 (
            .O(N__25617),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_));
    CascadeMux I__3773 (
            .O(N__25614),
            .I(N__25610));
    CascadeMux I__3772 (
            .O(N__25613),
            .I(N__25607));
    InMux I__3771 (
            .O(N__25610),
            .I(N__25602));
    InMux I__3770 (
            .O(N__25607),
            .I(N__25602));
    LocalMux I__3769 (
            .O(N__25602),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    InMux I__3768 (
            .O(N__25599),
            .I(N__25596));
    LocalMux I__3767 (
            .O(N__25596),
            .I(N__25593));
    Odrv4 I__3766 (
            .O(N__25593),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    InMux I__3765 (
            .O(N__25590),
            .I(N__25587));
    LocalMux I__3764 (
            .O(N__25587),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    CascadeMux I__3763 (
            .O(N__25584),
            .I(N__25581));
    InMux I__3762 (
            .O(N__25581),
            .I(N__25578));
    LocalMux I__3761 (
            .O(N__25578),
            .I(N__25575));
    Odrv4 I__3760 (
            .O(N__25575),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__3759 (
            .O(N__25572),
            .I(N__25569));
    LocalMux I__3758 (
            .O(N__25569),
            .I(N__25566));
    Odrv4 I__3757 (
            .O(N__25566),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    CascadeMux I__3756 (
            .O(N__25563),
            .I(N__25560));
    InMux I__3755 (
            .O(N__25560),
            .I(N__25557));
    LocalMux I__3754 (
            .O(N__25557),
            .I(N__25554));
    Odrv4 I__3753 (
            .O(N__25554),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    CascadeMux I__3752 (
            .O(N__25551),
            .I(N__25548));
    InMux I__3751 (
            .O(N__25548),
            .I(N__25545));
    LocalMux I__3750 (
            .O(N__25545),
            .I(N__25542));
    Span12Mux_s5_v I__3749 (
            .O(N__25542),
            .I(N__25539));
    Odrv12 I__3748 (
            .O(N__25539),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    InMux I__3747 (
            .O(N__25536),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__3746 (
            .O(N__25533),
            .I(N__25530));
    InMux I__3745 (
            .O(N__25530),
            .I(N__25527));
    LocalMux I__3744 (
            .O(N__25527),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    CascadeMux I__3743 (
            .O(N__25524),
            .I(N__25521));
    InMux I__3742 (
            .O(N__25521),
            .I(N__25518));
    LocalMux I__3741 (
            .O(N__25518),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__3740 (
            .O(N__25515),
            .I(N__25512));
    InMux I__3739 (
            .O(N__25512),
            .I(N__25509));
    LocalMux I__3738 (
            .O(N__25509),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__3737 (
            .O(N__25506),
            .I(N__25503));
    LocalMux I__3736 (
            .O(N__25503),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__3735 (
            .O(N__25500),
            .I(N__25497));
    InMux I__3734 (
            .O(N__25497),
            .I(N__25494));
    LocalMux I__3733 (
            .O(N__25494),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__3732 (
            .O(N__25491),
            .I(N__25488));
    InMux I__3731 (
            .O(N__25488),
            .I(N__25485));
    LocalMux I__3730 (
            .O(N__25485),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__3729 (
            .O(N__25482),
            .I(N__25479));
    InMux I__3728 (
            .O(N__25479),
            .I(N__25476));
    LocalMux I__3727 (
            .O(N__25476),
            .I(N__25473));
    Odrv4 I__3726 (
            .O(N__25473),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__3725 (
            .O(N__25470),
            .I(N__25467));
    InMux I__3724 (
            .O(N__25467),
            .I(N__25464));
    LocalMux I__3723 (
            .O(N__25464),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__3722 (
            .O(N__25461),
            .I(N__25458));
    InMux I__3721 (
            .O(N__25458),
            .I(N__25455));
    LocalMux I__3720 (
            .O(N__25455),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__3719 (
            .O(N__25452),
            .I(N__25449));
    LocalMux I__3718 (
            .O(N__25449),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__3717 (
            .O(N__25446),
            .I(\pwm_generator_inst.counter_cry_8 ));
    CascadeMux I__3716 (
            .O(N__25443),
            .I(N__25440));
    InMux I__3715 (
            .O(N__25440),
            .I(N__25437));
    LocalMux I__3714 (
            .O(N__25437),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__3713 (
            .O(N__25434),
            .I(N__25431));
    LocalMux I__3712 (
            .O(N__25431),
            .I(N__25428));
    Span4Mux_s1_v I__3711 (
            .O(N__25428),
            .I(N__25425));
    Odrv4 I__3710 (
            .O(N__25425),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__3709 (
            .O(N__25422),
            .I(N__25419));
    InMux I__3708 (
            .O(N__25419),
            .I(N__25416));
    LocalMux I__3707 (
            .O(N__25416),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__3706 (
            .O(N__25413),
            .I(N__25410));
    InMux I__3705 (
            .O(N__25410),
            .I(N__25407));
    LocalMux I__3704 (
            .O(N__25407),
            .I(N__25404));
    Odrv4 I__3703 (
            .O(N__25404),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__3702 (
            .O(N__25401),
            .I(N__25398));
    InMux I__3701 (
            .O(N__25398),
            .I(N__25395));
    LocalMux I__3700 (
            .O(N__25395),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__3699 (
            .O(N__25392),
            .I(N__25389));
    LocalMux I__3698 (
            .O(N__25389),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__3697 (
            .O(N__25386),
            .I(N__25383));
    InMux I__3696 (
            .O(N__25383),
            .I(N__25380));
    LocalMux I__3695 (
            .O(N__25380),
            .I(N__25377));
    Odrv4 I__3694 (
            .O(N__25377),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__3693 (
            .O(N__25374),
            .I(N__25371));
    InMux I__3692 (
            .O(N__25371),
            .I(N__25368));
    LocalMux I__3691 (
            .O(N__25368),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__3690 (
            .O(N__25365),
            .I(N__25362));
    LocalMux I__3689 (
            .O(N__25362),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__3688 (
            .O(N__25359),
            .I(N__25356));
    InMux I__3687 (
            .O(N__25356),
            .I(N__25353));
    LocalMux I__3686 (
            .O(N__25353),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__3685 (
            .O(N__25350),
            .I(N__25347));
    InMux I__3684 (
            .O(N__25347),
            .I(N__25344));
    LocalMux I__3683 (
            .O(N__25344),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__3682 (
            .O(N__25341),
            .I(bfn_7_26_0_));
    InMux I__3681 (
            .O(N__25338),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__3680 (
            .O(N__25335),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__3679 (
            .O(N__25332),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__3678 (
            .O(N__25329),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__3677 (
            .O(N__25326),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__3676 (
            .O(N__25323),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__3675 (
            .O(N__25320),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__3674 (
            .O(N__25317),
            .I(bfn_7_27_0_));
    InMux I__3673 (
            .O(N__25314),
            .I(N__25308));
    InMux I__3672 (
            .O(N__25313),
            .I(N__25301));
    InMux I__3671 (
            .O(N__25312),
            .I(N__25301));
    InMux I__3670 (
            .O(N__25311),
            .I(N__25301));
    LocalMux I__3669 (
            .O(N__25308),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__3668 (
            .O(N__25301),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    CascadeMux I__3667 (
            .O(N__25296),
            .I(N__25293));
    InMux I__3666 (
            .O(N__25293),
            .I(N__25286));
    InMux I__3665 (
            .O(N__25292),
            .I(N__25286));
    InMux I__3664 (
            .O(N__25291),
            .I(N__25283));
    LocalMux I__3663 (
            .O(N__25286),
            .I(N__25280));
    LocalMux I__3662 (
            .O(N__25283),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__3661 (
            .O(N__25280),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__3660 (
            .O(N__25275),
            .I(N__25269));
    InMux I__3659 (
            .O(N__25274),
            .I(N__25266));
    InMux I__3658 (
            .O(N__25273),
            .I(N__25263));
    InMux I__3657 (
            .O(N__25272),
            .I(N__25260));
    LocalMux I__3656 (
            .O(N__25269),
            .I(N__25255));
    LocalMux I__3655 (
            .O(N__25266),
            .I(N__25255));
    LocalMux I__3654 (
            .O(N__25263),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__3653 (
            .O(N__25260),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__3652 (
            .O(N__25255),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__3651 (
            .O(N__25248),
            .I(N__25242));
    ClkMux I__3650 (
            .O(N__25247),
            .I(N__25242));
    GlobalMux I__3649 (
            .O(N__25242),
            .I(N__25239));
    gio2CtrlBuf I__3648 (
            .O(N__25239),
            .I(delay_tr_input_c_g));
    InMux I__3647 (
            .O(N__25236),
            .I(N__25233));
    LocalMux I__3646 (
            .O(N__25233),
            .I(N__25230));
    Odrv12 I__3645 (
            .O(N__25230),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ));
    InMux I__3644 (
            .O(N__25227),
            .I(N__25224));
    LocalMux I__3643 (
            .O(N__25224),
            .I(N__25221));
    Odrv12 I__3642 (
            .O(N__25221),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ));
    InMux I__3641 (
            .O(N__25218),
            .I(N__25215));
    LocalMux I__3640 (
            .O(N__25215),
            .I(N__25212));
    Odrv12 I__3639 (
            .O(N__25212),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ));
    CascadeMux I__3638 (
            .O(N__25209),
            .I(N__25206));
    InMux I__3637 (
            .O(N__25206),
            .I(N__25203));
    LocalMux I__3636 (
            .O(N__25203),
            .I(N__25200));
    Odrv12 I__3635 (
            .O(N__25200),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ));
    InMux I__3634 (
            .O(N__25197),
            .I(N__25194));
    LocalMux I__3633 (
            .O(N__25194),
            .I(N__25191));
    Odrv12 I__3632 (
            .O(N__25191),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ));
    InMux I__3631 (
            .O(N__25188),
            .I(N__25185));
    LocalMux I__3630 (
            .O(N__25185),
            .I(N__25182));
    Odrv12 I__3629 (
            .O(N__25182),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ));
    InMux I__3628 (
            .O(N__25179),
            .I(bfn_7_16_0_));
    InMux I__3627 (
            .O(N__25176),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__3626 (
            .O(N__25173),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__3625 (
            .O(N__25170),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__3624 (
            .O(N__25167),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__3623 (
            .O(N__25164),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__3622 (
            .O(N__25161),
            .I(N__25156));
    CEMux I__3621 (
            .O(N__25160),
            .I(N__25153));
    CEMux I__3620 (
            .O(N__25159),
            .I(N__25150));
    LocalMux I__3619 (
            .O(N__25156),
            .I(N__25146));
    LocalMux I__3618 (
            .O(N__25153),
            .I(N__25141));
    LocalMux I__3617 (
            .O(N__25150),
            .I(N__25141));
    CEMux I__3616 (
            .O(N__25149),
            .I(N__25138));
    Span4Mux_h I__3615 (
            .O(N__25146),
            .I(N__25135));
    Span4Mux_v I__3614 (
            .O(N__25141),
            .I(N__25132));
    LocalMux I__3613 (
            .O(N__25138),
            .I(N__25129));
    Odrv4 I__3612 (
            .O(N__25135),
            .I(\delay_measurement_inst.delay_tr_timer.N_166_i ));
    Odrv4 I__3611 (
            .O(N__25132),
            .I(\delay_measurement_inst.delay_tr_timer.N_166_i ));
    Odrv12 I__3610 (
            .O(N__25129),
            .I(\delay_measurement_inst.delay_tr_timer.N_166_i ));
    InMux I__3609 (
            .O(N__25122),
            .I(N__25084));
    InMux I__3608 (
            .O(N__25121),
            .I(N__25084));
    InMux I__3607 (
            .O(N__25120),
            .I(N__25084));
    InMux I__3606 (
            .O(N__25119),
            .I(N__25084));
    InMux I__3605 (
            .O(N__25118),
            .I(N__25075));
    InMux I__3604 (
            .O(N__25117),
            .I(N__25075));
    InMux I__3603 (
            .O(N__25116),
            .I(N__25075));
    InMux I__3602 (
            .O(N__25115),
            .I(N__25075));
    InMux I__3601 (
            .O(N__25114),
            .I(N__25066));
    InMux I__3600 (
            .O(N__25113),
            .I(N__25066));
    InMux I__3599 (
            .O(N__25112),
            .I(N__25066));
    InMux I__3598 (
            .O(N__25111),
            .I(N__25066));
    InMux I__3597 (
            .O(N__25110),
            .I(N__25057));
    InMux I__3596 (
            .O(N__25109),
            .I(N__25057));
    InMux I__3595 (
            .O(N__25108),
            .I(N__25057));
    InMux I__3594 (
            .O(N__25107),
            .I(N__25057));
    InMux I__3593 (
            .O(N__25106),
            .I(N__25048));
    InMux I__3592 (
            .O(N__25105),
            .I(N__25048));
    InMux I__3591 (
            .O(N__25104),
            .I(N__25048));
    InMux I__3590 (
            .O(N__25103),
            .I(N__25048));
    InMux I__3589 (
            .O(N__25102),
            .I(N__25039));
    InMux I__3588 (
            .O(N__25101),
            .I(N__25039));
    InMux I__3587 (
            .O(N__25100),
            .I(N__25039));
    InMux I__3586 (
            .O(N__25099),
            .I(N__25039));
    InMux I__3585 (
            .O(N__25098),
            .I(N__25034));
    InMux I__3584 (
            .O(N__25097),
            .I(N__25034));
    InMux I__3583 (
            .O(N__25096),
            .I(N__25025));
    InMux I__3582 (
            .O(N__25095),
            .I(N__25025));
    InMux I__3581 (
            .O(N__25094),
            .I(N__25025));
    InMux I__3580 (
            .O(N__25093),
            .I(N__25025));
    LocalMux I__3579 (
            .O(N__25084),
            .I(N__25012));
    LocalMux I__3578 (
            .O(N__25075),
            .I(N__25012));
    LocalMux I__3577 (
            .O(N__25066),
            .I(N__25012));
    LocalMux I__3576 (
            .O(N__25057),
            .I(N__25012));
    LocalMux I__3575 (
            .O(N__25048),
            .I(N__25012));
    LocalMux I__3574 (
            .O(N__25039),
            .I(N__25012));
    LocalMux I__3573 (
            .O(N__25034),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__3572 (
            .O(N__25025),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv12 I__3571 (
            .O(N__25012),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__3570 (
            .O(N__25005),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__3569 (
            .O(N__25002),
            .I(bfn_7_15_0_));
    InMux I__3568 (
            .O(N__24999),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__3567 (
            .O(N__24996),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__3566 (
            .O(N__24993),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__3565 (
            .O(N__24990),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__3564 (
            .O(N__24987),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__3563 (
            .O(N__24984),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__3562 (
            .O(N__24981),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__3561 (
            .O(N__24978),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__3560 (
            .O(N__24975),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__3559 (
            .O(N__24972),
            .I(bfn_7_14_0_));
    InMux I__3558 (
            .O(N__24969),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__3557 (
            .O(N__24966),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__3556 (
            .O(N__24963),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__3555 (
            .O(N__24960),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__3554 (
            .O(N__24957),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__3553 (
            .O(N__24954),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__3552 (
            .O(N__24951),
            .I(bfn_7_13_0_));
    InMux I__3551 (
            .O(N__24948),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__3550 (
            .O(N__24945),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__3549 (
            .O(N__24942),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__3548 (
            .O(N__24939),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__3547 (
            .O(N__24936),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__3546 (
            .O(N__24933),
            .I(N__24927));
    InMux I__3545 (
            .O(N__24932),
            .I(N__24927));
    LocalMux I__3544 (
            .O(N__24927),
            .I(N__24924));
    Odrv4 I__3543 (
            .O(N__24924),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    InMux I__3542 (
            .O(N__24921),
            .I(N__24918));
    LocalMux I__3541 (
            .O(N__24918),
            .I(N__24914));
    InMux I__3540 (
            .O(N__24917),
            .I(N__24910));
    Span4Mux_v I__3539 (
            .O(N__24914),
            .I(N__24907));
    InMux I__3538 (
            .O(N__24913),
            .I(N__24904));
    LocalMux I__3537 (
            .O(N__24910),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv4 I__3536 (
            .O(N__24907),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    LocalMux I__3535 (
            .O(N__24904),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__3534 (
            .O(N__24897),
            .I(N__24892));
    InMux I__3533 (
            .O(N__24896),
            .I(N__24889));
    InMux I__3532 (
            .O(N__24895),
            .I(N__24886));
    LocalMux I__3531 (
            .O(N__24892),
            .I(N__24883));
    LocalMux I__3530 (
            .O(N__24889),
            .I(N__24880));
    LocalMux I__3529 (
            .O(N__24886),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    Odrv12 I__3528 (
            .O(N__24883),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    Odrv4 I__3527 (
            .O(N__24880),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    InMux I__3526 (
            .O(N__24873),
            .I(N__24867));
    InMux I__3525 (
            .O(N__24872),
            .I(N__24867));
    LocalMux I__3524 (
            .O(N__24867),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    CascadeMux I__3523 (
            .O(N__24864),
            .I(N__24860));
    InMux I__3522 (
            .O(N__24863),
            .I(N__24855));
    InMux I__3521 (
            .O(N__24860),
            .I(N__24855));
    LocalMux I__3520 (
            .O(N__24855),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    InMux I__3519 (
            .O(N__24852),
            .I(N__24849));
    LocalMux I__3518 (
            .O(N__24849),
            .I(N__24844));
    InMux I__3517 (
            .O(N__24848),
            .I(N__24841));
    InMux I__3516 (
            .O(N__24847),
            .I(N__24838));
    Span4Mux_h I__3515 (
            .O(N__24844),
            .I(N__24835));
    LocalMux I__3514 (
            .O(N__24841),
            .I(N__24832));
    LocalMux I__3513 (
            .O(N__24838),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv4 I__3512 (
            .O(N__24835),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv4 I__3511 (
            .O(N__24832),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    InMux I__3510 (
            .O(N__24825),
            .I(N__24821));
    InMux I__3509 (
            .O(N__24824),
            .I(N__24818));
    LocalMux I__3508 (
            .O(N__24821),
            .I(N__24813));
    LocalMux I__3507 (
            .O(N__24818),
            .I(N__24813));
    Odrv4 I__3506 (
            .O(N__24813),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__3505 (
            .O(N__24810),
            .I(N__24806));
    CascadeMux I__3504 (
            .O(N__24809),
            .I(N__24803));
    InMux I__3503 (
            .O(N__24806),
            .I(N__24800));
    InMux I__3502 (
            .O(N__24803),
            .I(N__24797));
    LocalMux I__3501 (
            .O(N__24800),
            .I(N__24792));
    LocalMux I__3500 (
            .O(N__24797),
            .I(N__24792));
    Odrv12 I__3499 (
            .O(N__24792),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__3498 (
            .O(N__24789),
            .I(N__24786));
    LocalMux I__3497 (
            .O(N__24786),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__3496 (
            .O(N__24783),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__3495 (
            .O(N__24780),
            .I(N__24777));
    LocalMux I__3494 (
            .O(N__24777),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__3493 (
            .O(N__24774),
            .I(bfn_5_25_0_));
    CascadeMux I__3492 (
            .O(N__24771),
            .I(N__24767));
    InMux I__3491 (
            .O(N__24770),
            .I(N__24761));
    InMux I__3490 (
            .O(N__24767),
            .I(N__24758));
    CascadeMux I__3489 (
            .O(N__24766),
            .I(N__24752));
    CascadeMux I__3488 (
            .O(N__24765),
            .I(N__24749));
    CascadeMux I__3487 (
            .O(N__24764),
            .I(N__24746));
    LocalMux I__3486 (
            .O(N__24761),
            .I(N__24742));
    LocalMux I__3485 (
            .O(N__24758),
            .I(N__24739));
    InMux I__3484 (
            .O(N__24757),
            .I(N__24733));
    InMux I__3483 (
            .O(N__24756),
            .I(N__24730));
    InMux I__3482 (
            .O(N__24755),
            .I(N__24721));
    InMux I__3481 (
            .O(N__24752),
            .I(N__24721));
    InMux I__3480 (
            .O(N__24749),
            .I(N__24721));
    InMux I__3479 (
            .O(N__24746),
            .I(N__24721));
    InMux I__3478 (
            .O(N__24745),
            .I(N__24718));
    Span4Mux_v I__3477 (
            .O(N__24742),
            .I(N__24713));
    Span4Mux_v I__3476 (
            .O(N__24739),
            .I(N__24713));
    InMux I__3475 (
            .O(N__24738),
            .I(N__24706));
    InMux I__3474 (
            .O(N__24737),
            .I(N__24706));
    InMux I__3473 (
            .O(N__24736),
            .I(N__24706));
    LocalMux I__3472 (
            .O(N__24733),
            .I(N__24697));
    LocalMux I__3471 (
            .O(N__24730),
            .I(N__24697));
    LocalMux I__3470 (
            .O(N__24721),
            .I(N__24697));
    LocalMux I__3469 (
            .O(N__24718),
            .I(N__24697));
    Odrv4 I__3468 (
            .O(N__24713),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    LocalMux I__3467 (
            .O(N__24706),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv12 I__3466 (
            .O(N__24697),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__3465 (
            .O(N__24690),
            .I(N__24687));
    LocalMux I__3464 (
            .O(N__24687),
            .I(N__24684));
    Span4Mux_h I__3463 (
            .O(N__24684),
            .I(N__24681));
    Span4Mux_h I__3462 (
            .O(N__24681),
            .I(N__24678));
    Odrv4 I__3461 (
            .O(N__24678),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    CascadeMux I__3460 (
            .O(N__24675),
            .I(N__24672));
    InMux I__3459 (
            .O(N__24672),
            .I(N__24669));
    LocalMux I__3458 (
            .O(N__24669),
            .I(N__24666));
    Span12Mux_h I__3457 (
            .O(N__24666),
            .I(N__24663));
    Odrv12 I__3456 (
            .O(N__24663),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    InMux I__3455 (
            .O(N__24660),
            .I(N__24657));
    LocalMux I__3454 (
            .O(N__24657),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__3453 (
            .O(N__24654),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__3452 (
            .O(N__24651),
            .I(N__24648));
    LocalMux I__3451 (
            .O(N__24648),
            .I(N__24645));
    Span4Mux_h I__3450 (
            .O(N__24645),
            .I(N__24642));
    Span4Mux_h I__3449 (
            .O(N__24642),
            .I(N__24639));
    Odrv4 I__3448 (
            .O(N__24639),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    CascadeMux I__3447 (
            .O(N__24636),
            .I(N__24633));
    InMux I__3446 (
            .O(N__24633),
            .I(N__24630));
    LocalMux I__3445 (
            .O(N__24630),
            .I(N__24627));
    Span4Mux_h I__3444 (
            .O(N__24627),
            .I(N__24624));
    Sp12to4 I__3443 (
            .O(N__24624),
            .I(N__24621));
    Span12Mux_h I__3442 (
            .O(N__24621),
            .I(N__24618));
    Odrv12 I__3441 (
            .O(N__24618),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    InMux I__3440 (
            .O(N__24615),
            .I(N__24612));
    LocalMux I__3439 (
            .O(N__24612),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__3438 (
            .O(N__24609),
            .I(bfn_5_24_0_));
    InMux I__3437 (
            .O(N__24606),
            .I(N__24603));
    LocalMux I__3436 (
            .O(N__24603),
            .I(N__24600));
    Span4Mux_h I__3435 (
            .O(N__24600),
            .I(N__24597));
    Span4Mux_h I__3434 (
            .O(N__24597),
            .I(N__24594));
    Odrv4 I__3433 (
            .O(N__24594),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    CascadeMux I__3432 (
            .O(N__24591),
            .I(N__24588));
    InMux I__3431 (
            .O(N__24588),
            .I(N__24585));
    LocalMux I__3430 (
            .O(N__24585),
            .I(N__24582));
    Span4Mux_h I__3429 (
            .O(N__24582),
            .I(N__24579));
    Sp12to4 I__3428 (
            .O(N__24579),
            .I(N__24576));
    Span12Mux_h I__3427 (
            .O(N__24576),
            .I(N__24573));
    Odrv12 I__3426 (
            .O(N__24573),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    InMux I__3425 (
            .O(N__24570),
            .I(N__24567));
    LocalMux I__3424 (
            .O(N__24567),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__3423 (
            .O(N__24564),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    CascadeMux I__3422 (
            .O(N__24561),
            .I(N__24558));
    InMux I__3421 (
            .O(N__24558),
            .I(N__24555));
    LocalMux I__3420 (
            .O(N__24555),
            .I(N__24552));
    Span4Mux_h I__3419 (
            .O(N__24552),
            .I(N__24549));
    Sp12to4 I__3418 (
            .O(N__24549),
            .I(N__24546));
    Span12Mux_h I__3417 (
            .O(N__24546),
            .I(N__24543));
    Odrv12 I__3416 (
            .O(N__24543),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__3415 (
            .O(N__24540),
            .I(N__24537));
    LocalMux I__3414 (
            .O(N__24537),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__3413 (
            .O(N__24534),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    InMux I__3412 (
            .O(N__24531),
            .I(N__24528));
    LocalMux I__3411 (
            .O(N__24528),
            .I(N__24525));
    Span12Mux_s6_h I__3410 (
            .O(N__24525),
            .I(N__24522));
    Span12Mux_h I__3409 (
            .O(N__24522),
            .I(N__24519));
    Odrv12 I__3408 (
            .O(N__24519),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__3407 (
            .O(N__24516),
            .I(N__24513));
    LocalMux I__3406 (
            .O(N__24513),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__3405 (
            .O(N__24510),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    CascadeMux I__3404 (
            .O(N__24507),
            .I(N__24504));
    InMux I__3403 (
            .O(N__24504),
            .I(N__24501));
    LocalMux I__3402 (
            .O(N__24501),
            .I(N__24498));
    Span12Mux_h I__3401 (
            .O(N__24498),
            .I(N__24495));
    Odrv12 I__3400 (
            .O(N__24495),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__3399 (
            .O(N__24492),
            .I(N__24489));
    LocalMux I__3398 (
            .O(N__24489),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__3397 (
            .O(N__24486),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    InMux I__3396 (
            .O(N__24483),
            .I(N__24480));
    LocalMux I__3395 (
            .O(N__24480),
            .I(N__24477));
    Span12Mux_h I__3394 (
            .O(N__24477),
            .I(N__24474));
    Odrv12 I__3393 (
            .O(N__24474),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__3392 (
            .O(N__24471),
            .I(N__24468));
    LocalMux I__3391 (
            .O(N__24468),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__3390 (
            .O(N__24465),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    CascadeMux I__3389 (
            .O(N__24462),
            .I(N__24459));
    InMux I__3388 (
            .O(N__24459),
            .I(N__24456));
    LocalMux I__3387 (
            .O(N__24456),
            .I(N__24453));
    Sp12to4 I__3386 (
            .O(N__24453),
            .I(N__24450));
    Span12Mux_s11_h I__3385 (
            .O(N__24450),
            .I(N__24447));
    Span12Mux_h I__3384 (
            .O(N__24447),
            .I(N__24444));
    Odrv12 I__3383 (
            .O(N__24444),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__3382 (
            .O(N__24441),
            .I(N__24438));
    LocalMux I__3381 (
            .O(N__24438),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__3380 (
            .O(N__24435),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    InMux I__3379 (
            .O(N__24432),
            .I(N__24429));
    LocalMux I__3378 (
            .O(N__24429),
            .I(N__24426));
    Span12Mux_s9_h I__3377 (
            .O(N__24426),
            .I(N__24423));
    Span12Mux_h I__3376 (
            .O(N__24423),
            .I(N__24420));
    Odrv12 I__3375 (
            .O(N__24420),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__3374 (
            .O(N__24417),
            .I(N__24414));
    InMux I__3373 (
            .O(N__24414),
            .I(N__24411));
    LocalMux I__3372 (
            .O(N__24411),
            .I(N__24408));
    Span4Mux_h I__3371 (
            .O(N__24408),
            .I(N__24405));
    Span4Mux_h I__3370 (
            .O(N__24405),
            .I(N__24402));
    Odrv4 I__3369 (
            .O(N__24402),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__3368 (
            .O(N__24399),
            .I(N__24396));
    LocalMux I__3367 (
            .O(N__24396),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__3366 (
            .O(N__24393),
            .I(N__24390));
    LocalMux I__3365 (
            .O(N__24390),
            .I(N__24387));
    Span4Mux_h I__3364 (
            .O(N__24387),
            .I(N__24384));
    Sp12to4 I__3363 (
            .O(N__24384),
            .I(N__24381));
    Span12Mux_h I__3362 (
            .O(N__24381),
            .I(N__24378));
    Odrv12 I__3361 (
            .O(N__24378),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__3360 (
            .O(N__24375),
            .I(N__24372));
    InMux I__3359 (
            .O(N__24372),
            .I(N__24369));
    LocalMux I__3358 (
            .O(N__24369),
            .I(N__24366));
    Span4Mux_h I__3357 (
            .O(N__24366),
            .I(N__24363));
    Span4Mux_h I__3356 (
            .O(N__24363),
            .I(N__24360));
    Odrv4 I__3355 (
            .O(N__24360),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    InMux I__3354 (
            .O(N__24357),
            .I(N__24354));
    LocalMux I__3353 (
            .O(N__24354),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__3352 (
            .O(N__24351),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__3351 (
            .O(N__24348),
            .I(N__24345));
    LocalMux I__3350 (
            .O(N__24345),
            .I(N__24342));
    Span12Mux_s7_h I__3349 (
            .O(N__24342),
            .I(N__24339));
    Span12Mux_h I__3348 (
            .O(N__24339),
            .I(N__24336));
    Odrv12 I__3347 (
            .O(N__24336),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__3346 (
            .O(N__24333),
            .I(N__24330));
    InMux I__3345 (
            .O(N__24330),
            .I(N__24327));
    LocalMux I__3344 (
            .O(N__24327),
            .I(N__24324));
    Span4Mux_h I__3343 (
            .O(N__24324),
            .I(N__24321));
    Span4Mux_h I__3342 (
            .O(N__24321),
            .I(N__24318));
    Odrv4 I__3341 (
            .O(N__24318),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    CascadeMux I__3340 (
            .O(N__24315),
            .I(N__24312));
    InMux I__3339 (
            .O(N__24312),
            .I(N__24309));
    LocalMux I__3338 (
            .O(N__24309),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__3337 (
            .O(N__24306),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__3336 (
            .O(N__24303),
            .I(N__24300));
    LocalMux I__3335 (
            .O(N__24300),
            .I(N__24297));
    Span12Mux_s6_h I__3334 (
            .O(N__24297),
            .I(N__24294));
    Span12Mux_h I__3333 (
            .O(N__24294),
            .I(N__24291));
    Odrv12 I__3332 (
            .O(N__24291),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__3331 (
            .O(N__24288),
            .I(N__24285));
    InMux I__3330 (
            .O(N__24285),
            .I(N__24282));
    LocalMux I__3329 (
            .O(N__24282),
            .I(N__24279));
    Span12Mux_h I__3328 (
            .O(N__24279),
            .I(N__24276));
    Odrv12 I__3327 (
            .O(N__24276),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    InMux I__3326 (
            .O(N__24273),
            .I(N__24270));
    LocalMux I__3325 (
            .O(N__24270),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__3324 (
            .O(N__24267),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__3323 (
            .O(N__24264),
            .I(N__24261));
    LocalMux I__3322 (
            .O(N__24261),
            .I(N__24258));
    Span12Mux_v I__3321 (
            .O(N__24258),
            .I(N__24255));
    Odrv12 I__3320 (
            .O(N__24255),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    CascadeMux I__3319 (
            .O(N__24252),
            .I(N__24249));
    InMux I__3318 (
            .O(N__24249),
            .I(N__24246));
    LocalMux I__3317 (
            .O(N__24246),
            .I(N__24243));
    Span12Mux_h I__3316 (
            .O(N__24243),
            .I(N__24240));
    Odrv12 I__3315 (
            .O(N__24240),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    InMux I__3314 (
            .O(N__24237),
            .I(N__24234));
    LocalMux I__3313 (
            .O(N__24234),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__3312 (
            .O(N__24231),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__3311 (
            .O(N__24228),
            .I(N__24225));
    LocalMux I__3310 (
            .O(N__24225),
            .I(N__24222));
    Span12Mux_h I__3309 (
            .O(N__24222),
            .I(N__24219));
    Odrv12 I__3308 (
            .O(N__24219),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__3307 (
            .O(N__24216),
            .I(N__24213));
    InMux I__3306 (
            .O(N__24213),
            .I(N__24210));
    LocalMux I__3305 (
            .O(N__24210),
            .I(N__24207));
    Span4Mux_h I__3304 (
            .O(N__24207),
            .I(N__24204));
    Span4Mux_h I__3303 (
            .O(N__24204),
            .I(N__24201));
    Odrv4 I__3302 (
            .O(N__24201),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__3301 (
            .O(N__24198),
            .I(N__24195));
    LocalMux I__3300 (
            .O(N__24195),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__3299 (
            .O(N__24192),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__3298 (
            .O(N__24189),
            .I(N__24186));
    LocalMux I__3297 (
            .O(N__24186),
            .I(N__24183));
    Span4Mux_h I__3296 (
            .O(N__24183),
            .I(N__24180));
    Span4Mux_h I__3295 (
            .O(N__24180),
            .I(N__24177));
    Odrv4 I__3294 (
            .O(N__24177),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    CascadeMux I__3293 (
            .O(N__24174),
            .I(N__24171));
    InMux I__3292 (
            .O(N__24171),
            .I(N__24168));
    LocalMux I__3291 (
            .O(N__24168),
            .I(N__24165));
    Span12Mux_h I__3290 (
            .O(N__24165),
            .I(N__24162));
    Odrv12 I__3289 (
            .O(N__24162),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    InMux I__3288 (
            .O(N__24159),
            .I(N__24156));
    LocalMux I__3287 (
            .O(N__24156),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__3286 (
            .O(N__24153),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__3285 (
            .O(N__24150),
            .I(N__24147));
    LocalMux I__3284 (
            .O(N__24147),
            .I(N__24143));
    InMux I__3283 (
            .O(N__24146),
            .I(N__24140));
    Odrv12 I__3282 (
            .O(N__24143),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    LocalMux I__3281 (
            .O(N__24140),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    CascadeMux I__3280 (
            .O(N__24135),
            .I(N__24132));
    InMux I__3279 (
            .O(N__24132),
            .I(N__24129));
    LocalMux I__3278 (
            .O(N__24129),
            .I(N__24126));
    Odrv4 I__3277 (
            .O(N__24126),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__3276 (
            .O(N__24123),
            .I(N__24118));
    InMux I__3275 (
            .O(N__24122),
            .I(N__24115));
    InMux I__3274 (
            .O(N__24121),
            .I(N__24112));
    LocalMux I__3273 (
            .O(N__24118),
            .I(N__24109));
    LocalMux I__3272 (
            .O(N__24115),
            .I(N__24106));
    LocalMux I__3271 (
            .O(N__24112),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__3270 (
            .O(N__24109),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__3269 (
            .O(N__24106),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__3268 (
            .O(N__24099),
            .I(N__24096));
    LocalMux I__3267 (
            .O(N__24096),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__3266 (
            .O(N__24093),
            .I(N__24089));
    InMux I__3265 (
            .O(N__24092),
            .I(N__24086));
    LocalMux I__3264 (
            .O(N__24089),
            .I(N__24083));
    LocalMux I__3263 (
            .O(N__24086),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    Odrv4 I__3262 (
            .O(N__24083),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    InMux I__3261 (
            .O(N__24078),
            .I(N__24075));
    LocalMux I__3260 (
            .O(N__24075),
            .I(N__24072));
    Odrv4 I__3259 (
            .O(N__24072),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    CascadeMux I__3258 (
            .O(N__24069),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ));
    CascadeMux I__3257 (
            .O(N__24066),
            .I(N__24062));
    InMux I__3256 (
            .O(N__24065),
            .I(N__24057));
    InMux I__3255 (
            .O(N__24062),
            .I(N__24057));
    LocalMux I__3254 (
            .O(N__24057),
            .I(N__24054));
    Odrv4 I__3253 (
            .O(N__24054),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__3252 (
            .O(N__24051),
            .I(N__24048));
    LocalMux I__3251 (
            .O(N__24048),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__3250 (
            .O(N__24045),
            .I(N__24042));
    LocalMux I__3249 (
            .O(N__24042),
            .I(N__24039));
    Span4Mux_v I__3248 (
            .O(N__24039),
            .I(N__24036));
    Odrv4 I__3247 (
            .O(N__24036),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    InMux I__3246 (
            .O(N__24033),
            .I(N__24030));
    LocalMux I__3245 (
            .O(N__24030),
            .I(N__24027));
    Span4Mux_v I__3244 (
            .O(N__24027),
            .I(N__24024));
    Span4Mux_h I__3243 (
            .O(N__24024),
            .I(N__24021));
    Odrv4 I__3242 (
            .O(N__24021),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ));
    InMux I__3241 (
            .O(N__24018),
            .I(N__24015));
    LocalMux I__3240 (
            .O(N__24015),
            .I(N__24012));
    Span4Mux_h I__3239 (
            .O(N__24012),
            .I(N__24009));
    Odrv4 I__3238 (
            .O(N__24009),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ));
    InMux I__3237 (
            .O(N__24006),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__3236 (
            .O(N__24003),
            .I(N__24000));
    LocalMux I__3235 (
            .O(N__24000),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ));
    InMux I__3234 (
            .O(N__23997),
            .I(N__23994));
    LocalMux I__3233 (
            .O(N__23994),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ));
    CascadeMux I__3232 (
            .O(N__23991),
            .I(N__23988));
    InMux I__3231 (
            .O(N__23988),
            .I(N__23985));
    LocalMux I__3230 (
            .O(N__23985),
            .I(N__23982));
    Odrv4 I__3229 (
            .O(N__23982),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ));
    InMux I__3228 (
            .O(N__23979),
            .I(N__23976));
    LocalMux I__3227 (
            .O(N__23976),
            .I(N__23973));
    Odrv4 I__3226 (
            .O(N__23973),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    CascadeMux I__3225 (
            .O(N__23970),
            .I(N__23967));
    InMux I__3224 (
            .O(N__23967),
            .I(N__23962));
    InMux I__3223 (
            .O(N__23966),
            .I(N__23959));
    InMux I__3222 (
            .O(N__23965),
            .I(N__23956));
    LocalMux I__3221 (
            .O(N__23962),
            .I(N__23953));
    LocalMux I__3220 (
            .O(N__23959),
            .I(N__23950));
    LocalMux I__3219 (
            .O(N__23956),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__3218 (
            .O(N__23953),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__3217 (
            .O(N__23950),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__3216 (
            .O(N__23943),
            .I(N__23940));
    LocalMux I__3215 (
            .O(N__23940),
            .I(N__23936));
    InMux I__3214 (
            .O(N__23939),
            .I(N__23933));
    Odrv12 I__3213 (
            .O(N__23936),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    LocalMux I__3212 (
            .O(N__23933),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__3211 (
            .O(N__23928),
            .I(N__23925));
    LocalMux I__3210 (
            .O(N__23925),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    InMux I__3209 (
            .O(N__23922),
            .I(N__23919));
    LocalMux I__3208 (
            .O(N__23919),
            .I(N__23916));
    Span4Mux_h I__3207 (
            .O(N__23916),
            .I(N__23912));
    InMux I__3206 (
            .O(N__23915),
            .I(N__23909));
    Odrv4 I__3205 (
            .O(N__23912),
            .I(\pwm_generator_inst.O_10 ));
    LocalMux I__3204 (
            .O(N__23909),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__3203 (
            .O(N__23904),
            .I(N__23901));
    LocalMux I__3202 (
            .O(N__23901),
            .I(N__23898));
    Span4Mux_v I__3201 (
            .O(N__23898),
            .I(N__23894));
    InMux I__3200 (
            .O(N__23897),
            .I(N__23890));
    Span4Mux_h I__3199 (
            .O(N__23894),
            .I(N__23887));
    InMux I__3198 (
            .O(N__23893),
            .I(N__23884));
    LocalMux I__3197 (
            .O(N__23890),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__3196 (
            .O(N__23887),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    LocalMux I__3195 (
            .O(N__23884),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    CascadeMux I__3194 (
            .O(N__23877),
            .I(N__23874));
    InMux I__3193 (
            .O(N__23874),
            .I(N__23871));
    LocalMux I__3192 (
            .O(N__23871),
            .I(N__23868));
    Odrv4 I__3191 (
            .O(N__23868),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    InMux I__3190 (
            .O(N__23865),
            .I(N__23862));
    LocalMux I__3189 (
            .O(N__23862),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    CascadeMux I__3188 (
            .O(N__23859),
            .I(N__23856));
    InMux I__3187 (
            .O(N__23856),
            .I(N__23853));
    LocalMux I__3186 (
            .O(N__23853),
            .I(N__23850));
    Span4Mux_h I__3185 (
            .O(N__23850),
            .I(N__23847));
    Odrv4 I__3184 (
            .O(N__23847),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    InMux I__3183 (
            .O(N__23844),
            .I(bfn_4_23_0_));
    InMux I__3182 (
            .O(N__23841),
            .I(N__23837));
    InMux I__3181 (
            .O(N__23840),
            .I(N__23834));
    LocalMux I__3180 (
            .O(N__23837),
            .I(N__23831));
    LocalMux I__3179 (
            .O(N__23834),
            .I(N__23828));
    Span4Mux_h I__3178 (
            .O(N__23831),
            .I(N__23825));
    Span4Mux_v I__3177 (
            .O(N__23828),
            .I(N__23822));
    Odrv4 I__3176 (
            .O(N__23825),
            .I(\pwm_generator_inst.un3_threshold ));
    Odrv4 I__3175 (
            .O(N__23822),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__3174 (
            .O(N__23817),
            .I(N__23814));
    LocalMux I__3173 (
            .O(N__23814),
            .I(N__23811));
    Span4Mux_h I__3172 (
            .O(N__23811),
            .I(N__23808));
    Odrv4 I__3171 (
            .O(N__23808),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__3170 (
            .O(N__23805),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__3169 (
            .O(N__23802),
            .I(N__23799));
    LocalMux I__3168 (
            .O(N__23799),
            .I(N__23796));
    Span4Mux_v I__3167 (
            .O(N__23796),
            .I(N__23793));
    Odrv4 I__3166 (
            .O(N__23793),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__3165 (
            .O(N__23790),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__3164 (
            .O(N__23787),
            .I(N__23784));
    LocalMux I__3163 (
            .O(N__23784),
            .I(N__23781));
    Span4Mux_h I__3162 (
            .O(N__23781),
            .I(N__23778));
    Odrv4 I__3161 (
            .O(N__23778),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__3160 (
            .O(N__23775),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__3159 (
            .O(N__23772),
            .I(N__23769));
    LocalMux I__3158 (
            .O(N__23769),
            .I(N__23766));
    Span4Mux_h I__3157 (
            .O(N__23766),
            .I(N__23762));
    InMux I__3156 (
            .O(N__23765),
            .I(N__23759));
    Odrv4 I__3155 (
            .O(N__23762),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    LocalMux I__3154 (
            .O(N__23759),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    InMux I__3153 (
            .O(N__23754),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    CascadeMux I__3152 (
            .O(N__23751),
            .I(N__23747));
    InMux I__3151 (
            .O(N__23750),
            .I(N__23742));
    InMux I__3150 (
            .O(N__23747),
            .I(N__23742));
    LocalMux I__3149 (
            .O(N__23742),
            .I(N__23739));
    Odrv4 I__3148 (
            .O(N__23739),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    InMux I__3147 (
            .O(N__23736),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__3146 (
            .O(N__23733),
            .I(N__23730));
    LocalMux I__3145 (
            .O(N__23730),
            .I(N__23726));
    InMux I__3144 (
            .O(N__23729),
            .I(N__23723));
    Odrv4 I__3143 (
            .O(N__23726),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    LocalMux I__3142 (
            .O(N__23723),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    InMux I__3141 (
            .O(N__23718),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__3140 (
            .O(N__23715),
            .I(N__23711));
    InMux I__3139 (
            .O(N__23714),
            .I(N__23708));
    LocalMux I__3138 (
            .O(N__23711),
            .I(N__23705));
    LocalMux I__3137 (
            .O(N__23708),
            .I(N__23702));
    Span4Mux_v I__3136 (
            .O(N__23705),
            .I(N__23699));
    Odrv4 I__3135 (
            .O(N__23702),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    Odrv4 I__3134 (
            .O(N__23699),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    InMux I__3133 (
            .O(N__23694),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    CascadeMux I__3132 (
            .O(N__23691),
            .I(N__23688));
    InMux I__3131 (
            .O(N__23688),
            .I(N__23685));
    LocalMux I__3130 (
            .O(N__23685),
            .I(N__23682));
    Odrv4 I__3129 (
            .O(N__23682),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    InMux I__3128 (
            .O(N__23679),
            .I(N__23676));
    LocalMux I__3127 (
            .O(N__23676),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__3126 (
            .O(N__23673),
            .I(N__23670));
    LocalMux I__3125 (
            .O(N__23670),
            .I(N__23667));
    Odrv4 I__3124 (
            .O(N__23667),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    InMux I__3123 (
            .O(N__23664),
            .I(N__23661));
    LocalMux I__3122 (
            .O(N__23661),
            .I(N__23658));
    Span4Mux_h I__3121 (
            .O(N__23658),
            .I(N__23655));
    Odrv4 I__3120 (
            .O(N__23655),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ));
    InMux I__3119 (
            .O(N__23652),
            .I(N__23649));
    LocalMux I__3118 (
            .O(N__23649),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    InMux I__3117 (
            .O(N__23646),
            .I(N__23643));
    LocalMux I__3116 (
            .O(N__23643),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ));
    InMux I__3115 (
            .O(N__23640),
            .I(N__23637));
    LocalMux I__3114 (
            .O(N__23637),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    CascadeMux I__3113 (
            .O(N__23634),
            .I(N__23631));
    InMux I__3112 (
            .O(N__23631),
            .I(N__23628));
    LocalMux I__3111 (
            .O(N__23628),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    InMux I__3110 (
            .O(N__23625),
            .I(N__23622));
    LocalMux I__3109 (
            .O(N__23622),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    InMux I__3108 (
            .O(N__23619),
            .I(N__23616));
    LocalMux I__3107 (
            .O(N__23616),
            .I(N__23613));
    Span4Mux_v I__3106 (
            .O(N__23613),
            .I(N__23610));
    Odrv4 I__3105 (
            .O(N__23610),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__3104 (
            .O(N__23607),
            .I(N__23604));
    LocalMux I__3103 (
            .O(N__23604),
            .I(N__23601));
    Odrv4 I__3102 (
            .O(N__23601),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__3101 (
            .O(N__23598),
            .I(N__23594));
    InMux I__3100 (
            .O(N__23597),
            .I(N__23575));
    LocalMux I__3099 (
            .O(N__23594),
            .I(N__23572));
    InMux I__3098 (
            .O(N__23593),
            .I(N__23567));
    InMux I__3097 (
            .O(N__23592),
            .I(N__23567));
    InMux I__3096 (
            .O(N__23591),
            .I(N__23564));
    InMux I__3095 (
            .O(N__23590),
            .I(N__23561));
    InMux I__3094 (
            .O(N__23589),
            .I(N__23556));
    InMux I__3093 (
            .O(N__23588),
            .I(N__23556));
    InMux I__3092 (
            .O(N__23587),
            .I(N__23553));
    InMux I__3091 (
            .O(N__23586),
            .I(N__23549));
    InMux I__3090 (
            .O(N__23585),
            .I(N__23534));
    InMux I__3089 (
            .O(N__23584),
            .I(N__23534));
    InMux I__3088 (
            .O(N__23583),
            .I(N__23534));
    InMux I__3087 (
            .O(N__23582),
            .I(N__23534));
    InMux I__3086 (
            .O(N__23581),
            .I(N__23534));
    InMux I__3085 (
            .O(N__23580),
            .I(N__23534));
    InMux I__3084 (
            .O(N__23579),
            .I(N__23534));
    InMux I__3083 (
            .O(N__23578),
            .I(N__23531));
    LocalMux I__3082 (
            .O(N__23575),
            .I(N__23510));
    Span4Mux_h I__3081 (
            .O(N__23572),
            .I(N__23510));
    LocalMux I__3080 (
            .O(N__23567),
            .I(N__23510));
    LocalMux I__3079 (
            .O(N__23564),
            .I(N__23510));
    LocalMux I__3078 (
            .O(N__23561),
            .I(N__23507));
    LocalMux I__3077 (
            .O(N__23556),
            .I(N__23501));
    LocalMux I__3076 (
            .O(N__23553),
            .I(N__23501));
    InMux I__3075 (
            .O(N__23552),
            .I(N__23498));
    LocalMux I__3074 (
            .O(N__23549),
            .I(N__23491));
    LocalMux I__3073 (
            .O(N__23534),
            .I(N__23491));
    LocalMux I__3072 (
            .O(N__23531),
            .I(N__23491));
    InMux I__3071 (
            .O(N__23530),
            .I(N__23488));
    InMux I__3070 (
            .O(N__23529),
            .I(N__23477));
    InMux I__3069 (
            .O(N__23528),
            .I(N__23477));
    InMux I__3068 (
            .O(N__23527),
            .I(N__23477));
    InMux I__3067 (
            .O(N__23526),
            .I(N__23477));
    InMux I__3066 (
            .O(N__23525),
            .I(N__23477));
    InMux I__3065 (
            .O(N__23524),
            .I(N__23474));
    InMux I__3064 (
            .O(N__23523),
            .I(N__23463));
    InMux I__3063 (
            .O(N__23522),
            .I(N__23463));
    InMux I__3062 (
            .O(N__23521),
            .I(N__23463));
    InMux I__3061 (
            .O(N__23520),
            .I(N__23463));
    InMux I__3060 (
            .O(N__23519),
            .I(N__23463));
    Span4Mux_v I__3059 (
            .O(N__23510),
            .I(N__23458));
    Span4Mux_v I__3058 (
            .O(N__23507),
            .I(N__23458));
    InMux I__3057 (
            .O(N__23506),
            .I(N__23455));
    Span4Mux_v I__3056 (
            .O(N__23501),
            .I(N__23450));
    LocalMux I__3055 (
            .O(N__23498),
            .I(N__23450));
    Span4Mux_v I__3054 (
            .O(N__23491),
            .I(N__23445));
    LocalMux I__3053 (
            .O(N__23488),
            .I(N__23445));
    LocalMux I__3052 (
            .O(N__23477),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3051 (
            .O(N__23474),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3050 (
            .O(N__23463),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3049 (
            .O(N__23458),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3048 (
            .O(N__23455),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3047 (
            .O(N__23450),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3046 (
            .O(N__23445),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__3045 (
            .O(N__23430),
            .I(N__23412));
    InMux I__3044 (
            .O(N__23429),
            .I(N__23412));
    InMux I__3043 (
            .O(N__23428),
            .I(N__23409));
    InMux I__3042 (
            .O(N__23427),
            .I(N__23406));
    InMux I__3041 (
            .O(N__23426),
            .I(N__23391));
    InMux I__3040 (
            .O(N__23425),
            .I(N__23391));
    InMux I__3039 (
            .O(N__23424),
            .I(N__23391));
    InMux I__3038 (
            .O(N__23423),
            .I(N__23391));
    InMux I__3037 (
            .O(N__23422),
            .I(N__23391));
    InMux I__3036 (
            .O(N__23421),
            .I(N__23391));
    InMux I__3035 (
            .O(N__23420),
            .I(N__23391));
    InMux I__3034 (
            .O(N__23419),
            .I(N__23382));
    InMux I__3033 (
            .O(N__23418),
            .I(N__23382));
    CascadeMux I__3032 (
            .O(N__23417),
            .I(N__23375));
    LocalMux I__3031 (
            .O(N__23412),
            .I(N__23366));
    LocalMux I__3030 (
            .O(N__23409),
            .I(N__23359));
    LocalMux I__3029 (
            .O(N__23406),
            .I(N__23359));
    LocalMux I__3028 (
            .O(N__23391),
            .I(N__23359));
    InMux I__3027 (
            .O(N__23390),
            .I(N__23352));
    InMux I__3026 (
            .O(N__23389),
            .I(N__23352));
    InMux I__3025 (
            .O(N__23388),
            .I(N__23352));
    InMux I__3024 (
            .O(N__23387),
            .I(N__23349));
    LocalMux I__3023 (
            .O(N__23382),
            .I(N__23346));
    InMux I__3022 (
            .O(N__23381),
            .I(N__23341));
    InMux I__3021 (
            .O(N__23380),
            .I(N__23341));
    CascadeMux I__3020 (
            .O(N__23379),
            .I(N__23335));
    CascadeMux I__3019 (
            .O(N__23378),
            .I(N__23332));
    InMux I__3018 (
            .O(N__23375),
            .I(N__23329));
    InMux I__3017 (
            .O(N__23374),
            .I(N__23318));
    InMux I__3016 (
            .O(N__23373),
            .I(N__23318));
    InMux I__3015 (
            .O(N__23372),
            .I(N__23318));
    InMux I__3014 (
            .O(N__23371),
            .I(N__23318));
    InMux I__3013 (
            .O(N__23370),
            .I(N__23318));
    InMux I__3012 (
            .O(N__23369),
            .I(N__23315));
    Span4Mux_h I__3011 (
            .O(N__23366),
            .I(N__23312));
    Span4Mux_h I__3010 (
            .O(N__23359),
            .I(N__23305));
    LocalMux I__3009 (
            .O(N__23352),
            .I(N__23305));
    LocalMux I__3008 (
            .O(N__23349),
            .I(N__23305));
    Span4Mux_h I__3007 (
            .O(N__23346),
            .I(N__23300));
    LocalMux I__3006 (
            .O(N__23341),
            .I(N__23300));
    InMux I__3005 (
            .O(N__23340),
            .I(N__23289));
    InMux I__3004 (
            .O(N__23339),
            .I(N__23289));
    InMux I__3003 (
            .O(N__23338),
            .I(N__23289));
    InMux I__3002 (
            .O(N__23335),
            .I(N__23289));
    InMux I__3001 (
            .O(N__23332),
            .I(N__23289));
    LocalMux I__3000 (
            .O(N__23329),
            .I(N__23284));
    LocalMux I__2999 (
            .O(N__23318),
            .I(N__23284));
    LocalMux I__2998 (
            .O(N__23315),
            .I(N__23279));
    Span4Mux_v I__2997 (
            .O(N__23312),
            .I(N__23279));
    Span4Mux_v I__2996 (
            .O(N__23305),
            .I(N__23276));
    Span4Mux_v I__2995 (
            .O(N__23300),
            .I(N__23273));
    LocalMux I__2994 (
            .O(N__23289),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2993 (
            .O(N__23284),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2992 (
            .O(N__23279),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2991 (
            .O(N__23276),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__2990 (
            .O(N__23273),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    CascadeMux I__2989 (
            .O(N__23262),
            .I(N__23259));
    InMux I__2988 (
            .O(N__23259),
            .I(N__23256));
    LocalMux I__2987 (
            .O(N__23256),
            .I(N__23253));
    Span4Mux_h I__2986 (
            .O(N__23253),
            .I(N__23250));
    Odrv4 I__2985 (
            .O(N__23250),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    CascadeMux I__2984 (
            .O(N__23247),
            .I(N__23234));
    CascadeMux I__2983 (
            .O(N__23246),
            .I(N__23231));
    CascadeMux I__2982 (
            .O(N__23245),
            .I(N__23227));
    CascadeMux I__2981 (
            .O(N__23244),
            .I(N__23224));
    CascadeMux I__2980 (
            .O(N__23243),
            .I(N__23218));
    CascadeMux I__2979 (
            .O(N__23242),
            .I(N__23214));
    CascadeMux I__2978 (
            .O(N__23241),
            .I(N__23209));
    CascadeMux I__2977 (
            .O(N__23240),
            .I(N__23197));
    CascadeMux I__2976 (
            .O(N__23239),
            .I(N__23193));
    CascadeMux I__2975 (
            .O(N__23238),
            .I(N__23190));
    CascadeMux I__2974 (
            .O(N__23237),
            .I(N__23187));
    InMux I__2973 (
            .O(N__23234),
            .I(N__23182));
    InMux I__2972 (
            .O(N__23231),
            .I(N__23182));
    InMux I__2971 (
            .O(N__23230),
            .I(N__23179));
    InMux I__2970 (
            .O(N__23227),
            .I(N__23172));
    InMux I__2969 (
            .O(N__23224),
            .I(N__23172));
    InMux I__2968 (
            .O(N__23223),
            .I(N__23172));
    InMux I__2967 (
            .O(N__23222),
            .I(N__23167));
    InMux I__2966 (
            .O(N__23221),
            .I(N__23167));
    InMux I__2965 (
            .O(N__23218),
            .I(N__23164));
    InMux I__2964 (
            .O(N__23217),
            .I(N__23159));
    InMux I__2963 (
            .O(N__23214),
            .I(N__23159));
    InMux I__2962 (
            .O(N__23213),
            .I(N__23152));
    InMux I__2961 (
            .O(N__23212),
            .I(N__23152));
    InMux I__2960 (
            .O(N__23209),
            .I(N__23152));
    CascadeMux I__2959 (
            .O(N__23208),
            .I(N__23146));
    CascadeMux I__2958 (
            .O(N__23207),
            .I(N__23143));
    CascadeMux I__2957 (
            .O(N__23206),
            .I(N__23140));
    InMux I__2956 (
            .O(N__23205),
            .I(N__23137));
    InMux I__2955 (
            .O(N__23204),
            .I(N__23126));
    InMux I__2954 (
            .O(N__23203),
            .I(N__23126));
    InMux I__2953 (
            .O(N__23202),
            .I(N__23126));
    InMux I__2952 (
            .O(N__23201),
            .I(N__23126));
    InMux I__2951 (
            .O(N__23200),
            .I(N__23126));
    InMux I__2950 (
            .O(N__23197),
            .I(N__23123));
    InMux I__2949 (
            .O(N__23196),
            .I(N__23114));
    InMux I__2948 (
            .O(N__23193),
            .I(N__23114));
    InMux I__2947 (
            .O(N__23190),
            .I(N__23114));
    InMux I__2946 (
            .O(N__23187),
            .I(N__23114));
    LocalMux I__2945 (
            .O(N__23182),
            .I(N__23111));
    LocalMux I__2944 (
            .O(N__23179),
            .I(N__23108));
    LocalMux I__2943 (
            .O(N__23172),
            .I(N__23105));
    LocalMux I__2942 (
            .O(N__23167),
            .I(N__23096));
    LocalMux I__2941 (
            .O(N__23164),
            .I(N__23096));
    LocalMux I__2940 (
            .O(N__23159),
            .I(N__23096));
    LocalMux I__2939 (
            .O(N__23152),
            .I(N__23096));
    InMux I__2938 (
            .O(N__23151),
            .I(N__23093));
    InMux I__2937 (
            .O(N__23150),
            .I(N__23082));
    InMux I__2936 (
            .O(N__23149),
            .I(N__23082));
    InMux I__2935 (
            .O(N__23146),
            .I(N__23082));
    InMux I__2934 (
            .O(N__23143),
            .I(N__23082));
    InMux I__2933 (
            .O(N__23140),
            .I(N__23082));
    LocalMux I__2932 (
            .O(N__23137),
            .I(N__23079));
    LocalMux I__2931 (
            .O(N__23126),
            .I(N__23076));
    LocalMux I__2930 (
            .O(N__23123),
            .I(N__23067));
    LocalMux I__2929 (
            .O(N__23114),
            .I(N__23067));
    Span4Mux_h I__2928 (
            .O(N__23111),
            .I(N__23067));
    Span4Mux_s3_h I__2927 (
            .O(N__23108),
            .I(N__23067));
    Span4Mux_s3_h I__2926 (
            .O(N__23105),
            .I(N__23062));
    Span4Mux_v I__2925 (
            .O(N__23096),
            .I(N__23062));
    LocalMux I__2924 (
            .O(N__23093),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    LocalMux I__2923 (
            .O(N__23082),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2922 (
            .O(N__23079),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2921 (
            .O(N__23076),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2920 (
            .O(N__23067),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2919 (
            .O(N__23062),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    InMux I__2918 (
            .O(N__23049),
            .I(N__23046));
    LocalMux I__2917 (
            .O(N__23046),
            .I(N__23043));
    Odrv4 I__2916 (
            .O(N__23043),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__2915 (
            .O(N__23040),
            .I(N__23037));
    LocalMux I__2914 (
            .O(N__23037),
            .I(N__23034));
    Span4Mux_v I__2913 (
            .O(N__23034),
            .I(N__23031));
    Odrv4 I__2912 (
            .O(N__23031),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__2911 (
            .O(N__23028),
            .I(N__23025));
    LocalMux I__2910 (
            .O(N__23025),
            .I(N__23022));
    Span4Mux_v I__2909 (
            .O(N__23022),
            .I(N__23019));
    Odrv4 I__2908 (
            .O(N__23019),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__2907 (
            .O(N__23016),
            .I(N__23013));
    InMux I__2906 (
            .O(N__23013),
            .I(N__23009));
    InMux I__2905 (
            .O(N__23012),
            .I(N__23004));
    LocalMux I__2904 (
            .O(N__23009),
            .I(N__23001));
    InMux I__2903 (
            .O(N__23008),
            .I(N__22998));
    InMux I__2902 (
            .O(N__23007),
            .I(N__22995));
    LocalMux I__2901 (
            .O(N__23004),
            .I(N__22992));
    Span4Mux_v I__2900 (
            .O(N__23001),
            .I(N__22987));
    LocalMux I__2899 (
            .O(N__22998),
            .I(N__22987));
    LocalMux I__2898 (
            .O(N__22995),
            .I(N__22984));
    Odrv4 I__2897 (
            .O(N__22992),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__2896 (
            .O(N__22987),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__2895 (
            .O(N__22984),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__2894 (
            .O(N__22977),
            .I(N__22974));
    InMux I__2893 (
            .O(N__22974),
            .I(N__22970));
    InMux I__2892 (
            .O(N__22973),
            .I(N__22966));
    LocalMux I__2891 (
            .O(N__22970),
            .I(N__22962));
    InMux I__2890 (
            .O(N__22969),
            .I(N__22959));
    LocalMux I__2889 (
            .O(N__22966),
            .I(N__22956));
    InMux I__2888 (
            .O(N__22965),
            .I(N__22953));
    Span4Mux_v I__2887 (
            .O(N__22962),
            .I(N__22946));
    LocalMux I__2886 (
            .O(N__22959),
            .I(N__22946));
    Span4Mux_h I__2885 (
            .O(N__22956),
            .I(N__22946));
    LocalMux I__2884 (
            .O(N__22953),
            .I(N__22943));
    Odrv4 I__2883 (
            .O(N__22946),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv12 I__2882 (
            .O(N__22943),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__2881 (
            .O(N__22938),
            .I(N__22935));
    InMux I__2880 (
            .O(N__22935),
            .I(N__22930));
    CascadeMux I__2879 (
            .O(N__22934),
            .I(N__22927));
    CascadeMux I__2878 (
            .O(N__22933),
            .I(N__22924));
    LocalMux I__2877 (
            .O(N__22930),
            .I(N__22921));
    InMux I__2876 (
            .O(N__22927),
            .I(N__22918));
    InMux I__2875 (
            .O(N__22924),
            .I(N__22914));
    Span12Mux_s3_h I__2874 (
            .O(N__22921),
            .I(N__22909));
    LocalMux I__2873 (
            .O(N__22918),
            .I(N__22909));
    InMux I__2872 (
            .O(N__22917),
            .I(N__22906));
    LocalMux I__2871 (
            .O(N__22914),
            .I(N__22903));
    Span12Mux_v I__2870 (
            .O(N__22909),
            .I(N__22900));
    LocalMux I__2869 (
            .O(N__22906),
            .I(N__22897));
    Odrv4 I__2868 (
            .O(N__22903),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv12 I__2867 (
            .O(N__22900),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__2866 (
            .O(N__22897),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__2865 (
            .O(N__22890),
            .I(N__22887));
    InMux I__2864 (
            .O(N__22887),
            .I(N__22884));
    LocalMux I__2863 (
            .O(N__22884),
            .I(N__22878));
    InMux I__2862 (
            .O(N__22883),
            .I(N__22875));
    InMux I__2861 (
            .O(N__22882),
            .I(N__22872));
    InMux I__2860 (
            .O(N__22881),
            .I(N__22869));
    Span4Mux_h I__2859 (
            .O(N__22878),
            .I(N__22864));
    LocalMux I__2858 (
            .O(N__22875),
            .I(N__22864));
    LocalMux I__2857 (
            .O(N__22872),
            .I(N__22861));
    LocalMux I__2856 (
            .O(N__22869),
            .I(N__22858));
    Span4Mux_v I__2855 (
            .O(N__22864),
            .I(N__22853));
    Span4Mux_v I__2854 (
            .O(N__22861),
            .I(N__22853));
    Odrv4 I__2853 (
            .O(N__22858),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__2852 (
            .O(N__22853),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__2851 (
            .O(N__22848),
            .I(N__22845));
    LocalMux I__2850 (
            .O(N__22845),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ));
    InMux I__2849 (
            .O(N__22842),
            .I(N__22839));
    LocalMux I__2848 (
            .O(N__22839),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__2847 (
            .O(N__22836),
            .I(N__22833));
    LocalMux I__2846 (
            .O(N__22833),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__2845 (
            .O(N__22830),
            .I(bfn_3_25_0_));
    InMux I__2844 (
            .O(N__22827),
            .I(N__22824));
    LocalMux I__2843 (
            .O(N__22824),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__2842 (
            .O(N__22821),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    InMux I__2841 (
            .O(N__22818),
            .I(N__22815));
    LocalMux I__2840 (
            .O(N__22815),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__2839 (
            .O(N__22812),
            .I(N__22805));
    InMux I__2838 (
            .O(N__22811),
            .I(N__22805));
    InMux I__2837 (
            .O(N__22810),
            .I(N__22802));
    LocalMux I__2836 (
            .O(N__22805),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__2835 (
            .O(N__22802),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__2834 (
            .O(N__22797),
            .I(N__22794));
    LocalMux I__2833 (
            .O(N__22794),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__2832 (
            .O(N__22791),
            .I(N__22788));
    LocalMux I__2831 (
            .O(N__22788),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    InMux I__2830 (
            .O(N__22785),
            .I(N__22780));
    InMux I__2829 (
            .O(N__22784),
            .I(N__22777));
    InMux I__2828 (
            .O(N__22783),
            .I(N__22774));
    LocalMux I__2827 (
            .O(N__22780),
            .I(N__22769));
    LocalMux I__2826 (
            .O(N__22777),
            .I(N__22769));
    LocalMux I__2825 (
            .O(N__22774),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv4 I__2824 (
            .O(N__22769),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__2823 (
            .O(N__22764),
            .I(N__22761));
    LocalMux I__2822 (
            .O(N__22761),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__2821 (
            .O(N__22758),
            .I(N__22751));
    InMux I__2820 (
            .O(N__22757),
            .I(N__22751));
    InMux I__2819 (
            .O(N__22756),
            .I(N__22748));
    LocalMux I__2818 (
            .O(N__22751),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__2817 (
            .O(N__22748),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    CascadeMux I__2816 (
            .O(N__22743),
            .I(N__22740));
    InMux I__2815 (
            .O(N__22740),
            .I(N__22737));
    LocalMux I__2814 (
            .O(N__22737),
            .I(N__22734));
    Odrv4 I__2813 (
            .O(N__22734),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__2812 (
            .O(N__22731),
            .I(N__22728));
    LocalMux I__2811 (
            .O(N__22728),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__2810 (
            .O(N__22725),
            .I(N__22722));
    LocalMux I__2809 (
            .O(N__22722),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__2808 (
            .O(N__22719),
            .I(N__22714));
    InMux I__2807 (
            .O(N__22718),
            .I(N__22711));
    InMux I__2806 (
            .O(N__22717),
            .I(N__22708));
    LocalMux I__2805 (
            .O(N__22714),
            .I(N__22705));
    LocalMux I__2804 (
            .O(N__22711),
            .I(N__22702));
    LocalMux I__2803 (
            .O(N__22708),
            .I(N__22697));
    Span4Mux_v I__2802 (
            .O(N__22705),
            .I(N__22697));
    Odrv4 I__2801 (
            .O(N__22702),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    Odrv4 I__2800 (
            .O(N__22697),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__2799 (
            .O(N__22692),
            .I(N__22689));
    LocalMux I__2798 (
            .O(N__22689),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    InMux I__2797 (
            .O(N__22686),
            .I(N__22683));
    LocalMux I__2796 (
            .O(N__22683),
            .I(N__22680));
    Span4Mux_v I__2795 (
            .O(N__22680),
            .I(N__22677));
    Span4Mux_h I__2794 (
            .O(N__22677),
            .I(N__22674));
    Odrv4 I__2793 (
            .O(N__22674),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    CascadeMux I__2792 (
            .O(N__22671),
            .I(N__22665));
    CascadeMux I__2791 (
            .O(N__22670),
            .I(N__22662));
    InMux I__2790 (
            .O(N__22669),
            .I(N__22659));
    InMux I__2789 (
            .O(N__22668),
            .I(N__22656));
    InMux I__2788 (
            .O(N__22665),
            .I(N__22653));
    InMux I__2787 (
            .O(N__22662),
            .I(N__22650));
    LocalMux I__2786 (
            .O(N__22659),
            .I(N__22643));
    LocalMux I__2785 (
            .O(N__22656),
            .I(N__22643));
    LocalMux I__2784 (
            .O(N__22653),
            .I(N__22643));
    LocalMux I__2783 (
            .O(N__22650),
            .I(N__22640));
    Span4Mux_v I__2782 (
            .O(N__22643),
            .I(N__22637));
    Span4Mux_v I__2781 (
            .O(N__22640),
            .I(N__22634));
    Odrv4 I__2780 (
            .O(N__22637),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__2779 (
            .O(N__22634),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__2778 (
            .O(N__22629),
            .I(N__22626));
    LocalMux I__2777 (
            .O(N__22626),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__2776 (
            .O(N__22623),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    InMux I__2775 (
            .O(N__22620),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__2774 (
            .O(N__22617),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__2773 (
            .O(N__22614),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__2772 (
            .O(N__22611),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__2771 (
            .O(N__22608),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__2770 (
            .O(N__22605),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    CascadeMux I__2769 (
            .O(N__22602),
            .I(N__22599));
    InMux I__2768 (
            .O(N__22599),
            .I(N__22596));
    LocalMux I__2767 (
            .O(N__22596),
            .I(N__22591));
    InMux I__2766 (
            .O(N__22595),
            .I(N__22587));
    InMux I__2765 (
            .O(N__22594),
            .I(N__22584));
    Span4Mux_v I__2764 (
            .O(N__22591),
            .I(N__22581));
    InMux I__2763 (
            .O(N__22590),
            .I(N__22578));
    LocalMux I__2762 (
            .O(N__22587),
            .I(N__22575));
    LocalMux I__2761 (
            .O(N__22584),
            .I(N__22572));
    Odrv4 I__2760 (
            .O(N__22581),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__2759 (
            .O(N__22578),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv12 I__2758 (
            .O(N__22575),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__2757 (
            .O(N__22572),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__2756 (
            .O(N__22563),
            .I(N__22559));
    CascadeMux I__2755 (
            .O(N__22562),
            .I(N__22556));
    InMux I__2754 (
            .O(N__22559),
            .I(N__22551));
    InMux I__2753 (
            .O(N__22556),
            .I(N__22551));
    LocalMux I__2752 (
            .O(N__22551),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2751 (
            .O(N__22548),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2750 (
            .O(N__22545),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2749 (
            .O(N__22542),
            .I(N__22539));
    LocalMux I__2748 (
            .O(N__22539),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    InMux I__2747 (
            .O(N__22536),
            .I(N__22533));
    LocalMux I__2746 (
            .O(N__22533),
            .I(N__22530));
    Odrv12 I__2745 (
            .O(N__22530),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__2744 (
            .O(N__22527),
            .I(N__22524));
    LocalMux I__2743 (
            .O(N__22524),
            .I(N__22521));
    Span4Mux_s3_h I__2742 (
            .O(N__22521),
            .I(N__22518));
    Odrv4 I__2741 (
            .O(N__22518),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    CascadeMux I__2740 (
            .O(N__22515),
            .I(N__22512));
    InMux I__2739 (
            .O(N__22512),
            .I(N__22508));
    InMux I__2738 (
            .O(N__22511),
            .I(N__22505));
    LocalMux I__2737 (
            .O(N__22508),
            .I(N__22501));
    LocalMux I__2736 (
            .O(N__22505),
            .I(N__22498));
    InMux I__2735 (
            .O(N__22504),
            .I(N__22495));
    Span12Mux_s3_h I__2734 (
            .O(N__22501),
            .I(N__22488));
    Sp12to4 I__2733 (
            .O(N__22498),
            .I(N__22488));
    LocalMux I__2732 (
            .O(N__22495),
            .I(N__22488));
    Odrv12 I__2731 (
            .O(N__22488),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2730 (
            .O(N__22485),
            .I(N__22481));
    InMux I__2729 (
            .O(N__22484),
            .I(N__22477));
    LocalMux I__2728 (
            .O(N__22481),
            .I(N__22474));
    InMux I__2727 (
            .O(N__22480),
            .I(N__22471));
    LocalMux I__2726 (
            .O(N__22477),
            .I(N__22468));
    Span4Mux_h I__2725 (
            .O(N__22474),
            .I(N__22463));
    LocalMux I__2724 (
            .O(N__22471),
            .I(N__22463));
    Span4Mux_v I__2723 (
            .O(N__22468),
            .I(N__22458));
    Span4Mux_v I__2722 (
            .O(N__22463),
            .I(N__22458));
    Odrv4 I__2721 (
            .O(N__22458),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    CascadeMux I__2720 (
            .O(N__22455),
            .I(N__22452));
    InMux I__2719 (
            .O(N__22452),
            .I(N__22449));
    LocalMux I__2718 (
            .O(N__22449),
            .I(N__22444));
    InMux I__2717 (
            .O(N__22448),
            .I(N__22441));
    InMux I__2716 (
            .O(N__22447),
            .I(N__22438));
    Span4Mux_v I__2715 (
            .O(N__22444),
            .I(N__22433));
    LocalMux I__2714 (
            .O(N__22441),
            .I(N__22433));
    LocalMux I__2713 (
            .O(N__22438),
            .I(N__22430));
    Span4Mux_v I__2712 (
            .O(N__22433),
            .I(N__22427));
    Odrv12 I__2711 (
            .O(N__22430),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2710 (
            .O(N__22427),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    CascadeMux I__2709 (
            .O(N__22422),
            .I(N__22419));
    InMux I__2708 (
            .O(N__22419),
            .I(N__22416));
    LocalMux I__2707 (
            .O(N__22416),
            .I(N__22411));
    InMux I__2706 (
            .O(N__22415),
            .I(N__22408));
    InMux I__2705 (
            .O(N__22414),
            .I(N__22405));
    Span4Mux_v I__2704 (
            .O(N__22411),
            .I(N__22400));
    LocalMux I__2703 (
            .O(N__22408),
            .I(N__22400));
    LocalMux I__2702 (
            .O(N__22405),
            .I(N__22397));
    Span4Mux_v I__2701 (
            .O(N__22400),
            .I(N__22394));
    Odrv12 I__2700 (
            .O(N__22397),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2699 (
            .O(N__22394),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    CascadeMux I__2698 (
            .O(N__22389),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    CascadeMux I__2697 (
            .O(N__22386),
            .I(N__22383));
    InMux I__2696 (
            .O(N__22383),
            .I(N__22379));
    InMux I__2695 (
            .O(N__22382),
            .I(N__22376));
    LocalMux I__2694 (
            .O(N__22379),
            .I(N__22372));
    LocalMux I__2693 (
            .O(N__22376),
            .I(N__22369));
    InMux I__2692 (
            .O(N__22375),
            .I(N__22366));
    Span4Mux_v I__2691 (
            .O(N__22372),
            .I(N__22363));
    Span4Mux_v I__2690 (
            .O(N__22369),
            .I(N__22358));
    LocalMux I__2689 (
            .O(N__22366),
            .I(N__22358));
    Span4Mux_v I__2688 (
            .O(N__22363),
            .I(N__22355));
    Span4Mux_v I__2687 (
            .O(N__22358),
            .I(N__22352));
    Odrv4 I__2686 (
            .O(N__22355),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__2685 (
            .O(N__22352),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    CascadeMux I__2684 (
            .O(N__22347),
            .I(N__22344));
    InMux I__2683 (
            .O(N__22344),
            .I(N__22341));
    LocalMux I__2682 (
            .O(N__22341),
            .I(N__22337));
    InMux I__2681 (
            .O(N__22340),
            .I(N__22334));
    Odrv4 I__2680 (
            .O(N__22337),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__2679 (
            .O(N__22334),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__2678 (
            .O(N__22329),
            .I(N__22326));
    LocalMux I__2677 (
            .O(N__22326),
            .I(N__22323));
    Odrv12 I__2676 (
            .O(N__22323),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__2675 (
            .O(N__22320),
            .I(N__22317));
    InMux I__2674 (
            .O(N__22317),
            .I(N__22312));
    CascadeMux I__2673 (
            .O(N__22316),
            .I(N__22309));
    CascadeMux I__2672 (
            .O(N__22315),
            .I(N__22306));
    LocalMux I__2671 (
            .O(N__22312),
            .I(N__22303));
    InMux I__2670 (
            .O(N__22309),
            .I(N__22299));
    InMux I__2669 (
            .O(N__22306),
            .I(N__22296));
    Span4Mux_v I__2668 (
            .O(N__22303),
            .I(N__22293));
    InMux I__2667 (
            .O(N__22302),
            .I(N__22290));
    LocalMux I__2666 (
            .O(N__22299),
            .I(N__22287));
    LocalMux I__2665 (
            .O(N__22296),
            .I(N__22284));
    Odrv4 I__2664 (
            .O(N__22293),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__2663 (
            .O(N__22290),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__2662 (
            .O(N__22287),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__2661 (
            .O(N__22284),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    CascadeMux I__2660 (
            .O(N__22275),
            .I(N__22272));
    InMux I__2659 (
            .O(N__22272),
            .I(N__22269));
    LocalMux I__2658 (
            .O(N__22269),
            .I(N__22266));
    Span4Mux_v I__2657 (
            .O(N__22266),
            .I(N__22262));
    InMux I__2656 (
            .O(N__22265),
            .I(N__22259));
    Odrv4 I__2655 (
            .O(N__22262),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    LocalMux I__2654 (
            .O(N__22259),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2653 (
            .O(N__22254),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__2652 (
            .O(N__22251),
            .I(N__22248));
    InMux I__2651 (
            .O(N__22248),
            .I(N__22244));
    CascadeMux I__2650 (
            .O(N__22247),
            .I(N__22241));
    LocalMux I__2649 (
            .O(N__22244),
            .I(N__22236));
    InMux I__2648 (
            .O(N__22241),
            .I(N__22233));
    InMux I__2647 (
            .O(N__22240),
            .I(N__22230));
    InMux I__2646 (
            .O(N__22239),
            .I(N__22227));
    Span4Mux_v I__2645 (
            .O(N__22236),
            .I(N__22224));
    LocalMux I__2644 (
            .O(N__22233),
            .I(N__22219));
    LocalMux I__2643 (
            .O(N__22230),
            .I(N__22219));
    LocalMux I__2642 (
            .O(N__22227),
            .I(N__22216));
    Odrv4 I__2641 (
            .O(N__22224),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__2640 (
            .O(N__22219),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv12 I__2639 (
            .O(N__22216),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__2638 (
            .O(N__22209),
            .I(N__22205));
    CascadeMux I__2637 (
            .O(N__22208),
            .I(N__22202));
    InMux I__2636 (
            .O(N__22205),
            .I(N__22197));
    InMux I__2635 (
            .O(N__22202),
            .I(N__22197));
    LocalMux I__2634 (
            .O(N__22197),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2633 (
            .O(N__22194),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2632 (
            .O(N__22191),
            .I(N__22187));
    CascadeMux I__2631 (
            .O(N__22190),
            .I(N__22183));
    LocalMux I__2630 (
            .O(N__22187),
            .I(N__22179));
    InMux I__2629 (
            .O(N__22186),
            .I(N__22176));
    InMux I__2628 (
            .O(N__22183),
            .I(N__22173));
    InMux I__2627 (
            .O(N__22182),
            .I(N__22170));
    Span4Mux_v I__2626 (
            .O(N__22179),
            .I(N__22165));
    LocalMux I__2625 (
            .O(N__22176),
            .I(N__22165));
    LocalMux I__2624 (
            .O(N__22173),
            .I(N__22162));
    LocalMux I__2623 (
            .O(N__22170),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__2622 (
            .O(N__22165),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__2621 (
            .O(N__22162),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__2620 (
            .O(N__22155),
            .I(N__22149));
    InMux I__2619 (
            .O(N__22154),
            .I(N__22149));
    LocalMux I__2618 (
            .O(N__22149),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2617 (
            .O(N__22146),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    CascadeMux I__2616 (
            .O(N__22143),
            .I(N__22140));
    InMux I__2615 (
            .O(N__22140),
            .I(N__22137));
    LocalMux I__2614 (
            .O(N__22137),
            .I(N__22132));
    CascadeMux I__2613 (
            .O(N__22136),
            .I(N__22129));
    InMux I__2612 (
            .O(N__22135),
            .I(N__22125));
    Span4Mux_v I__2611 (
            .O(N__22132),
            .I(N__22122));
    InMux I__2610 (
            .O(N__22129),
            .I(N__22119));
    InMux I__2609 (
            .O(N__22128),
            .I(N__22116));
    LocalMux I__2608 (
            .O(N__22125),
            .I(N__22113));
    Odrv4 I__2607 (
            .O(N__22122),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__2606 (
            .O(N__22119),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__2605 (
            .O(N__22116),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv12 I__2604 (
            .O(N__22113),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__2603 (
            .O(N__22104),
            .I(N__22101));
    LocalMux I__2602 (
            .O(N__22101),
            .I(N__22097));
    InMux I__2601 (
            .O(N__22100),
            .I(N__22094));
    Odrv4 I__2600 (
            .O(N__22097),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    LocalMux I__2599 (
            .O(N__22094),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2598 (
            .O(N__22089),
            .I(bfn_3_20_0_));
    CascadeMux I__2597 (
            .O(N__22086),
            .I(N__22083));
    InMux I__2596 (
            .O(N__22083),
            .I(N__22080));
    LocalMux I__2595 (
            .O(N__22080),
            .I(N__22077));
    Span4Mux_v I__2594 (
            .O(N__22077),
            .I(N__22072));
    InMux I__2593 (
            .O(N__22076),
            .I(N__22069));
    InMux I__2592 (
            .O(N__22075),
            .I(N__22065));
    Sp12to4 I__2591 (
            .O(N__22072),
            .I(N__22060));
    LocalMux I__2590 (
            .O(N__22069),
            .I(N__22060));
    InMux I__2589 (
            .O(N__22068),
            .I(N__22057));
    LocalMux I__2588 (
            .O(N__22065),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv12 I__2587 (
            .O(N__22060),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__2586 (
            .O(N__22057),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__2585 (
            .O(N__22050),
            .I(N__22046));
    CascadeMux I__2584 (
            .O(N__22049),
            .I(N__22043));
    LocalMux I__2583 (
            .O(N__22046),
            .I(N__22040));
    InMux I__2582 (
            .O(N__22043),
            .I(N__22037));
    Odrv4 I__2581 (
            .O(N__22040),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    LocalMux I__2580 (
            .O(N__22037),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2579 (
            .O(N__22032),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    CascadeMux I__2578 (
            .O(N__22029),
            .I(N__22026));
    InMux I__2577 (
            .O(N__22026),
            .I(N__22023));
    LocalMux I__2576 (
            .O(N__22023),
            .I(N__22020));
    Span4Mux_h I__2575 (
            .O(N__22020),
            .I(N__22014));
    InMux I__2574 (
            .O(N__22019),
            .I(N__22011));
    InMux I__2573 (
            .O(N__22018),
            .I(N__22008));
    InMux I__2572 (
            .O(N__22017),
            .I(N__22005));
    Span4Mux_v I__2571 (
            .O(N__22014),
            .I(N__22000));
    LocalMux I__2570 (
            .O(N__22011),
            .I(N__22000));
    LocalMux I__2569 (
            .O(N__22008),
            .I(N__21997));
    LocalMux I__2568 (
            .O(N__22005),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__2567 (
            .O(N__22000),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__2566 (
            .O(N__21997),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__2565 (
            .O(N__21990),
            .I(N__21984));
    InMux I__2564 (
            .O(N__21989),
            .I(N__21984));
    LocalMux I__2563 (
            .O(N__21984),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2562 (
            .O(N__21981),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    CascadeMux I__2561 (
            .O(N__21978),
            .I(N__21975));
    InMux I__2560 (
            .O(N__21975),
            .I(N__21971));
    CascadeMux I__2559 (
            .O(N__21974),
            .I(N__21967));
    LocalMux I__2558 (
            .O(N__21971),
            .I(N__21964));
    CascadeMux I__2557 (
            .O(N__21970),
            .I(N__21960));
    InMux I__2556 (
            .O(N__21967),
            .I(N__21957));
    Span4Mux_v I__2555 (
            .O(N__21964),
            .I(N__21954));
    InMux I__2554 (
            .O(N__21963),
            .I(N__21951));
    InMux I__2553 (
            .O(N__21960),
            .I(N__21948));
    LocalMux I__2552 (
            .O(N__21957),
            .I(N__21945));
    Odrv4 I__2551 (
            .O(N__21954),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__2550 (
            .O(N__21951),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__2549 (
            .O(N__21948),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv12 I__2548 (
            .O(N__21945),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__2547 (
            .O(N__21936),
            .I(N__21932));
    InMux I__2546 (
            .O(N__21935),
            .I(N__21929));
    LocalMux I__2545 (
            .O(N__21932),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__2544 (
            .O(N__21929),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2543 (
            .O(N__21924),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    CascadeMux I__2542 (
            .O(N__21921),
            .I(N__21918));
    InMux I__2541 (
            .O(N__21918),
            .I(N__21915));
    LocalMux I__2540 (
            .O(N__21915),
            .I(N__21912));
    Span4Mux_h I__2539 (
            .O(N__21912),
            .I(N__21909));
    Span4Mux_v I__2538 (
            .O(N__21909),
            .I(N__21903));
    InMux I__2537 (
            .O(N__21908),
            .I(N__21900));
    InMux I__2536 (
            .O(N__21907),
            .I(N__21895));
    InMux I__2535 (
            .O(N__21906),
            .I(N__21895));
    Odrv4 I__2534 (
            .O(N__21903),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__2533 (
            .O(N__21900),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__2532 (
            .O(N__21895),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__2531 (
            .O(N__21888),
            .I(N__21882));
    InMux I__2530 (
            .O(N__21887),
            .I(N__21882));
    LocalMux I__2529 (
            .O(N__21882),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2528 (
            .O(N__21879),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__2527 (
            .O(N__21876),
            .I(N__21873));
    InMux I__2526 (
            .O(N__21873),
            .I(N__21869));
    InMux I__2525 (
            .O(N__21872),
            .I(N__21865));
    LocalMux I__2524 (
            .O(N__21869),
            .I(N__21862));
    InMux I__2523 (
            .O(N__21868),
            .I(N__21859));
    LocalMux I__2522 (
            .O(N__21865),
            .I(N__21853));
    Span4Mux_v I__2521 (
            .O(N__21862),
            .I(N__21853));
    LocalMux I__2520 (
            .O(N__21859),
            .I(N__21850));
    InMux I__2519 (
            .O(N__21858),
            .I(N__21847));
    Odrv4 I__2518 (
            .O(N__21853),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__2517 (
            .O(N__21850),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__2516 (
            .O(N__21847),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__2515 (
            .O(N__21840),
            .I(N__21834));
    InMux I__2514 (
            .O(N__21839),
            .I(N__21834));
    LocalMux I__2513 (
            .O(N__21834),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2512 (
            .O(N__21831),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2511 (
            .O(N__21828),
            .I(N__21825));
    LocalMux I__2510 (
            .O(N__21825),
            .I(N__21822));
    Span4Mux_s3_h I__2509 (
            .O(N__21822),
            .I(N__21818));
    InMux I__2508 (
            .O(N__21821),
            .I(N__21815));
    Odrv4 I__2507 (
            .O(N__21818),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2506 (
            .O(N__21815),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2505 (
            .O(N__21810),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__2504 (
            .O(N__21807),
            .I(N__21804));
    LocalMux I__2503 (
            .O(N__21804),
            .I(N__21801));
    Span4Mux_s3_h I__2502 (
            .O(N__21801),
            .I(N__21797));
    InMux I__2501 (
            .O(N__21800),
            .I(N__21794));
    Odrv4 I__2500 (
            .O(N__21797),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__2499 (
            .O(N__21794),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2498 (
            .O(N__21789),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    CascadeMux I__2497 (
            .O(N__21786),
            .I(N__21783));
    InMux I__2496 (
            .O(N__21783),
            .I(N__21780));
    LocalMux I__2495 (
            .O(N__21780),
            .I(N__21775));
    InMux I__2494 (
            .O(N__21779),
            .I(N__21771));
    InMux I__2493 (
            .O(N__21778),
            .I(N__21768));
    Span4Mux_v I__2492 (
            .O(N__21775),
            .I(N__21765));
    InMux I__2491 (
            .O(N__21774),
            .I(N__21762));
    LocalMux I__2490 (
            .O(N__21771),
            .I(N__21757));
    LocalMux I__2489 (
            .O(N__21768),
            .I(N__21757));
    Odrv4 I__2488 (
            .O(N__21765),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__2487 (
            .O(N__21762),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv12 I__2486 (
            .O(N__21757),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__2485 (
            .O(N__21750),
            .I(N__21744));
    InMux I__2484 (
            .O(N__21749),
            .I(N__21744));
    LocalMux I__2483 (
            .O(N__21744),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2482 (
            .O(N__21741),
            .I(bfn_3_19_0_));
    InMux I__2481 (
            .O(N__21738),
            .I(N__21735));
    LocalMux I__2480 (
            .O(N__21735),
            .I(N__21732));
    Span4Mux_v I__2479 (
            .O(N__21732),
            .I(N__21729));
    Odrv4 I__2478 (
            .O(N__21729),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    CascadeMux I__2477 (
            .O(N__21726),
            .I(N__21723));
    InMux I__2476 (
            .O(N__21723),
            .I(N__21720));
    LocalMux I__2475 (
            .O(N__21720),
            .I(N__21714));
    InMux I__2474 (
            .O(N__21719),
            .I(N__21711));
    InMux I__2473 (
            .O(N__21718),
            .I(N__21708));
    InMux I__2472 (
            .O(N__21717),
            .I(N__21705));
    Span4Mux_v I__2471 (
            .O(N__21714),
            .I(N__21700));
    LocalMux I__2470 (
            .O(N__21711),
            .I(N__21700));
    LocalMux I__2469 (
            .O(N__21708),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__2468 (
            .O(N__21705),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__2467 (
            .O(N__21700),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__2466 (
            .O(N__21693),
            .I(N__21689));
    InMux I__2465 (
            .O(N__21692),
            .I(N__21686));
    LocalMux I__2464 (
            .O(N__21689),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__2463 (
            .O(N__21686),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2462 (
            .O(N__21681),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    CascadeMux I__2461 (
            .O(N__21678),
            .I(N__21675));
    InMux I__2460 (
            .O(N__21675),
            .I(N__21671));
    InMux I__2459 (
            .O(N__21674),
            .I(N__21667));
    LocalMux I__2458 (
            .O(N__21671),
            .I(N__21664));
    InMux I__2457 (
            .O(N__21670),
            .I(N__21660));
    LocalMux I__2456 (
            .O(N__21667),
            .I(N__21657));
    Span4Mux_v I__2455 (
            .O(N__21664),
            .I(N__21654));
    InMux I__2454 (
            .O(N__21663),
            .I(N__21651));
    LocalMux I__2453 (
            .O(N__21660),
            .I(N__21646));
    Span4Mux_v I__2452 (
            .O(N__21657),
            .I(N__21646));
    Odrv4 I__2451 (
            .O(N__21654),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__2450 (
            .O(N__21651),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__2449 (
            .O(N__21646),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__2448 (
            .O(N__21639),
            .I(N__21635));
    InMux I__2447 (
            .O(N__21638),
            .I(N__21632));
    LocalMux I__2446 (
            .O(N__21635),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    LocalMux I__2445 (
            .O(N__21632),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2444 (
            .O(N__21627),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2443 (
            .O(N__21624),
            .I(N__21621));
    LocalMux I__2442 (
            .O(N__21621),
            .I(N__21615));
    InMux I__2441 (
            .O(N__21620),
            .I(N__21612));
    CascadeMux I__2440 (
            .O(N__21619),
            .I(N__21609));
    InMux I__2439 (
            .O(N__21618),
            .I(N__21606));
    Span4Mux_v I__2438 (
            .O(N__21615),
            .I(N__21601));
    LocalMux I__2437 (
            .O(N__21612),
            .I(N__21601));
    InMux I__2436 (
            .O(N__21609),
            .I(N__21598));
    LocalMux I__2435 (
            .O(N__21606),
            .I(N__21595));
    Odrv4 I__2434 (
            .O(N__21601),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__2433 (
            .O(N__21598),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv12 I__2432 (
            .O(N__21595),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__2431 (
            .O(N__21588),
            .I(N__21585));
    InMux I__2430 (
            .O(N__21585),
            .I(N__21581));
    InMux I__2429 (
            .O(N__21584),
            .I(N__21578));
    LocalMux I__2428 (
            .O(N__21581),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    LocalMux I__2427 (
            .O(N__21578),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2426 (
            .O(N__21573),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__2425 (
            .O(N__21570),
            .I(N__21567));
    InMux I__2424 (
            .O(N__21567),
            .I(N__21563));
    CascadeMux I__2423 (
            .O(N__21566),
            .I(N__21560));
    LocalMux I__2422 (
            .O(N__21563),
            .I(N__21555));
    InMux I__2421 (
            .O(N__21560),
            .I(N__21552));
    InMux I__2420 (
            .O(N__21559),
            .I(N__21549));
    InMux I__2419 (
            .O(N__21558),
            .I(N__21546));
    Span4Mux_v I__2418 (
            .O(N__21555),
            .I(N__21541));
    LocalMux I__2417 (
            .O(N__21552),
            .I(N__21541));
    LocalMux I__2416 (
            .O(N__21549),
            .I(N__21538));
    LocalMux I__2415 (
            .O(N__21546),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__2414 (
            .O(N__21541),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__2413 (
            .O(N__21538),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__2412 (
            .O(N__21531),
            .I(N__21525));
    InMux I__2411 (
            .O(N__21530),
            .I(N__21525));
    LocalMux I__2410 (
            .O(N__21525),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2409 (
            .O(N__21522),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2408 (
            .O(N__21519),
            .I(N__21516));
    LocalMux I__2407 (
            .O(N__21516),
            .I(N__21513));
    Odrv12 I__2406 (
            .O(N__21513),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__2405 (
            .O(N__21510),
            .I(N__21505));
    InMux I__2404 (
            .O(N__21509),
            .I(N__21502));
    InMux I__2403 (
            .O(N__21508),
            .I(N__21499));
    InMux I__2402 (
            .O(N__21505),
            .I(N__21496));
    LocalMux I__2401 (
            .O(N__21502),
            .I(N__21492));
    LocalMux I__2400 (
            .O(N__21499),
            .I(N__21487));
    LocalMux I__2399 (
            .O(N__21496),
            .I(N__21487));
    InMux I__2398 (
            .O(N__21495),
            .I(N__21484));
    Span4Mux_s3_h I__2397 (
            .O(N__21492),
            .I(N__21481));
    Odrv4 I__2396 (
            .O(N__21487),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__2395 (
            .O(N__21484),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__2394 (
            .O(N__21481),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__2393 (
            .O(N__21474),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    CascadeMux I__2392 (
            .O(N__21471),
            .I(N__21466));
    CascadeMux I__2391 (
            .O(N__21470),
            .I(N__21463));
    InMux I__2390 (
            .O(N__21469),
            .I(N__21460));
    InMux I__2389 (
            .O(N__21466),
            .I(N__21457));
    InMux I__2388 (
            .O(N__21463),
            .I(N__21454));
    LocalMux I__2387 (
            .O(N__21460),
            .I(N__21446));
    LocalMux I__2386 (
            .O(N__21457),
            .I(N__21446));
    LocalMux I__2385 (
            .O(N__21454),
            .I(N__21446));
    InMux I__2384 (
            .O(N__21453),
            .I(N__21443));
    Span4Mux_v I__2383 (
            .O(N__21446),
            .I(N__21440));
    LocalMux I__2382 (
            .O(N__21443),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__2381 (
            .O(N__21440),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__2380 (
            .O(N__21435),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2379 (
            .O(N__21432),
            .I(N__21427));
    CascadeMux I__2378 (
            .O(N__21431),
            .I(N__21424));
    InMux I__2377 (
            .O(N__21430),
            .I(N__21420));
    LocalMux I__2376 (
            .O(N__21427),
            .I(N__21417));
    InMux I__2375 (
            .O(N__21424),
            .I(N__21414));
    InMux I__2374 (
            .O(N__21423),
            .I(N__21411));
    LocalMux I__2373 (
            .O(N__21420),
            .I(N__21408));
    Sp12to4 I__2372 (
            .O(N__21417),
            .I(N__21401));
    LocalMux I__2371 (
            .O(N__21414),
            .I(N__21401));
    LocalMux I__2370 (
            .O(N__21411),
            .I(N__21401));
    Odrv4 I__2369 (
            .O(N__21408),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv12 I__2368 (
            .O(N__21401),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__2367 (
            .O(N__21396),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    InMux I__2366 (
            .O(N__21393),
            .I(N__21390));
    LocalMux I__2365 (
            .O(N__21390),
            .I(N__21387));
    Odrv12 I__2364 (
            .O(N__21387),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__2363 (
            .O(N__21384),
            .I(N__21381));
    InMux I__2362 (
            .O(N__21381),
            .I(N__21377));
    InMux I__2361 (
            .O(N__21380),
            .I(N__21373));
    LocalMux I__2360 (
            .O(N__21377),
            .I(N__21370));
    InMux I__2359 (
            .O(N__21376),
            .I(N__21367));
    LocalMux I__2358 (
            .O(N__21373),
            .I(N__21361));
    Span4Mux_h I__2357 (
            .O(N__21370),
            .I(N__21361));
    LocalMux I__2356 (
            .O(N__21367),
            .I(N__21358));
    InMux I__2355 (
            .O(N__21366),
            .I(N__21355));
    Span4Mux_v I__2354 (
            .O(N__21361),
            .I(N__21350));
    Span4Mux_v I__2353 (
            .O(N__21358),
            .I(N__21350));
    LocalMux I__2352 (
            .O(N__21355),
            .I(N__21347));
    Odrv4 I__2351 (
            .O(N__21350),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__2350 (
            .O(N__21347),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__2349 (
            .O(N__21342),
            .I(bfn_3_18_0_));
    InMux I__2348 (
            .O(N__21339),
            .I(N__21336));
    LocalMux I__2347 (
            .O(N__21336),
            .I(N__21333));
    Odrv12 I__2346 (
            .O(N__21333),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__2345 (
            .O(N__21330),
            .I(N__21326));
    InMux I__2344 (
            .O(N__21329),
            .I(N__21321));
    InMux I__2343 (
            .O(N__21326),
            .I(N__21321));
    LocalMux I__2342 (
            .O(N__21321),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2341 (
            .O(N__21318),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    CascadeMux I__2340 (
            .O(N__21315),
            .I(N__21312));
    InMux I__2339 (
            .O(N__21312),
            .I(N__21308));
    InMux I__2338 (
            .O(N__21311),
            .I(N__21303));
    LocalMux I__2337 (
            .O(N__21308),
            .I(N__21300));
    InMux I__2336 (
            .O(N__21307),
            .I(N__21297));
    InMux I__2335 (
            .O(N__21306),
            .I(N__21294));
    LocalMux I__2334 (
            .O(N__21303),
            .I(N__21289));
    Span4Mux_h I__2333 (
            .O(N__21300),
            .I(N__21289));
    LocalMux I__2332 (
            .O(N__21297),
            .I(N__21286));
    LocalMux I__2331 (
            .O(N__21294),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__2330 (
            .O(N__21289),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__2329 (
            .O(N__21286),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__2328 (
            .O(N__21279),
            .I(N__21273));
    InMux I__2327 (
            .O(N__21278),
            .I(N__21273));
    LocalMux I__2326 (
            .O(N__21273),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2325 (
            .O(N__21270),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2324 (
            .O(N__21267),
            .I(N__21264));
    LocalMux I__2323 (
            .O(N__21264),
            .I(N__21261));
    Odrv4 I__2322 (
            .O(N__21261),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    CascadeMux I__2321 (
            .O(N__21258),
            .I(N__21254));
    InMux I__2320 (
            .O(N__21257),
            .I(N__21250));
    InMux I__2319 (
            .O(N__21254),
            .I(N__21246));
    InMux I__2318 (
            .O(N__21253),
            .I(N__21243));
    LocalMux I__2317 (
            .O(N__21250),
            .I(N__21240));
    CascadeMux I__2316 (
            .O(N__21249),
            .I(N__21237));
    LocalMux I__2315 (
            .O(N__21246),
            .I(N__21234));
    LocalMux I__2314 (
            .O(N__21243),
            .I(N__21231));
    Span4Mux_h I__2313 (
            .O(N__21240),
            .I(N__21228));
    InMux I__2312 (
            .O(N__21237),
            .I(N__21225));
    Span4Mux_h I__2311 (
            .O(N__21234),
            .I(N__21222));
    Span4Mux_s2_h I__2310 (
            .O(N__21231),
            .I(N__21219));
    Odrv4 I__2309 (
            .O(N__21228),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__2308 (
            .O(N__21225),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__2307 (
            .O(N__21222),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__2306 (
            .O(N__21219),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__2305 (
            .O(N__21210),
            .I(N__21206));
    InMux I__2304 (
            .O(N__21209),
            .I(N__21203));
    LocalMux I__2303 (
            .O(N__21206),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2302 (
            .O(N__21203),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2301 (
            .O(N__21198),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2300 (
            .O(N__21195),
            .I(N__21189));
    InMux I__2299 (
            .O(N__21194),
            .I(N__21189));
    LocalMux I__2298 (
            .O(N__21189),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2297 (
            .O(N__21186),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__2296 (
            .O(N__21183),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ));
    InMux I__2295 (
            .O(N__21180),
            .I(N__21177));
    LocalMux I__2294 (
            .O(N__21177),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__2293 (
            .O(N__21174),
            .I(N__21171));
    LocalMux I__2292 (
            .O(N__21171),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    CascadeMux I__2291 (
            .O(N__21168),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ));
    InMux I__2290 (
            .O(N__21165),
            .I(N__21162));
    LocalMux I__2289 (
            .O(N__21162),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    InMux I__2288 (
            .O(N__21159),
            .I(N__21156));
    LocalMux I__2287 (
            .O(N__21156),
            .I(N__21152));
    InMux I__2286 (
            .O(N__21155),
            .I(N__21149));
    Span4Mux_h I__2285 (
            .O(N__21152),
            .I(N__21146));
    LocalMux I__2284 (
            .O(N__21149),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    Odrv4 I__2283 (
            .O(N__21146),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__2282 (
            .O(N__21141),
            .I(N__21138));
    InMux I__2281 (
            .O(N__21138),
            .I(N__21133));
    InMux I__2280 (
            .O(N__21137),
            .I(N__21130));
    InMux I__2279 (
            .O(N__21136),
            .I(N__21127));
    LocalMux I__2278 (
            .O(N__21133),
            .I(N__21124));
    LocalMux I__2277 (
            .O(N__21130),
            .I(N__21120));
    LocalMux I__2276 (
            .O(N__21127),
            .I(N__21117));
    Span4Mux_v I__2275 (
            .O(N__21124),
            .I(N__21114));
    InMux I__2274 (
            .O(N__21123),
            .I(N__21110));
    Span4Mux_v I__2273 (
            .O(N__21120),
            .I(N__21107));
    Span4Mux_v I__2272 (
            .O(N__21117),
            .I(N__21104));
    Span4Mux_s3_h I__2271 (
            .O(N__21114),
            .I(N__21101));
    InMux I__2270 (
            .O(N__21113),
            .I(N__21098));
    LocalMux I__2269 (
            .O(N__21110),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__2268 (
            .O(N__21107),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__2267 (
            .O(N__21104),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__2266 (
            .O(N__21101),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__2265 (
            .O(N__21098),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__2264 (
            .O(N__21087),
            .I(N__21084));
    LocalMux I__2263 (
            .O(N__21084),
            .I(N__21081));
    Span4Mux_v I__2262 (
            .O(N__21081),
            .I(N__21078));
    Odrv4 I__2261 (
            .O(N__21078),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__2260 (
            .O(N__21075),
            .I(N__21071));
    CascadeMux I__2259 (
            .O(N__21074),
            .I(N__21068));
    InMux I__2258 (
            .O(N__21071),
            .I(N__21064));
    InMux I__2257 (
            .O(N__21068),
            .I(N__21061));
    InMux I__2256 (
            .O(N__21067),
            .I(N__21058));
    LocalMux I__2255 (
            .O(N__21064),
            .I(N__21053));
    LocalMux I__2254 (
            .O(N__21061),
            .I(N__21053));
    LocalMux I__2253 (
            .O(N__21058),
            .I(N__21050));
    Span4Mux_v I__2252 (
            .O(N__21053),
            .I(N__21047));
    Span4Mux_s2_h I__2251 (
            .O(N__21050),
            .I(N__21044));
    Odrv4 I__2250 (
            .O(N__21047),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__2249 (
            .O(N__21044),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__2248 (
            .O(N__21039),
            .I(N__21036));
    LocalMux I__2247 (
            .O(N__21036),
            .I(N__21033));
    Span4Mux_h I__2246 (
            .O(N__21033),
            .I(N__21030));
    Span4Mux_v I__2245 (
            .O(N__21030),
            .I(N__21027));
    Odrv4 I__2244 (
            .O(N__21027),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2243 (
            .O(N__21024),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2242 (
            .O(N__21021),
            .I(N__21018));
    LocalMux I__2241 (
            .O(N__21018),
            .I(N__21013));
    InMux I__2240 (
            .O(N__21017),
            .I(N__21007));
    InMux I__2239 (
            .O(N__21016),
            .I(N__21007));
    Span4Mux_v I__2238 (
            .O(N__21013),
            .I(N__21004));
    InMux I__2237 (
            .O(N__21012),
            .I(N__21001));
    LocalMux I__2236 (
            .O(N__21007),
            .I(N__20998));
    Odrv4 I__2235 (
            .O(N__21004),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__2234 (
            .O(N__21001),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv12 I__2233 (
            .O(N__20998),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    CascadeMux I__2232 (
            .O(N__20991),
            .I(N__20988));
    InMux I__2231 (
            .O(N__20988),
            .I(N__20985));
    LocalMux I__2230 (
            .O(N__20985),
            .I(N__20982));
    Odrv12 I__2229 (
            .O(N__20982),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__2228 (
            .O(N__20979),
            .I(N__20976));
    LocalMux I__2227 (
            .O(N__20976),
            .I(N__20971));
    InMux I__2226 (
            .O(N__20975),
            .I(N__20968));
    InMux I__2225 (
            .O(N__20974),
            .I(N__20965));
    Span4Mux_s3_h I__2224 (
            .O(N__20971),
            .I(N__20962));
    LocalMux I__2223 (
            .O(N__20968),
            .I(N__20957));
    LocalMux I__2222 (
            .O(N__20965),
            .I(N__20957));
    Span4Mux_v I__2221 (
            .O(N__20962),
            .I(N__20954));
    Span4Mux_v I__2220 (
            .O(N__20957),
            .I(N__20951));
    Odrv4 I__2219 (
            .O(N__20954),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__2218 (
            .O(N__20951),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2217 (
            .O(N__20946),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2216 (
            .O(N__20943),
            .I(N__20940));
    LocalMux I__2215 (
            .O(N__20940),
            .I(N__20937));
    Odrv4 I__2214 (
            .O(N__20937),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2213 (
            .O(N__20934),
            .I(N__20931));
    InMux I__2212 (
            .O(N__20931),
            .I(N__20925));
    CascadeMux I__2211 (
            .O(N__20930),
            .I(N__20922));
    InMux I__2210 (
            .O(N__20929),
            .I(N__20917));
    InMux I__2209 (
            .O(N__20928),
            .I(N__20917));
    LocalMux I__2208 (
            .O(N__20925),
            .I(N__20914));
    InMux I__2207 (
            .O(N__20922),
            .I(N__20911));
    LocalMux I__2206 (
            .O(N__20917),
            .I(N__20908));
    Span4Mux_v I__2205 (
            .O(N__20914),
            .I(N__20905));
    LocalMux I__2204 (
            .O(N__20911),
            .I(N__20902));
    Odrv4 I__2203 (
            .O(N__20908),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__2202 (
            .O(N__20905),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__2201 (
            .O(N__20902),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__2200 (
            .O(N__20895),
            .I(N__20891));
    CascadeMux I__2199 (
            .O(N__20894),
            .I(N__20886));
    LocalMux I__2198 (
            .O(N__20891),
            .I(N__20883));
    InMux I__2197 (
            .O(N__20890),
            .I(N__20880));
    InMux I__2196 (
            .O(N__20889),
            .I(N__20875));
    InMux I__2195 (
            .O(N__20886),
            .I(N__20875));
    Span4Mux_s3_h I__2194 (
            .O(N__20883),
            .I(N__20872));
    LocalMux I__2193 (
            .O(N__20880),
            .I(N__20867));
    LocalMux I__2192 (
            .O(N__20875),
            .I(N__20867));
    Span4Mux_v I__2191 (
            .O(N__20872),
            .I(N__20864));
    Span4Mux_v I__2190 (
            .O(N__20867),
            .I(N__20861));
    Odrv4 I__2189 (
            .O(N__20864),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2188 (
            .O(N__20861),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2187 (
            .O(N__20856),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2186 (
            .O(N__20853),
            .I(N__20850));
    LocalMux I__2185 (
            .O(N__20850),
            .I(N__20847));
    Span4Mux_v I__2184 (
            .O(N__20847),
            .I(N__20844));
    Odrv4 I__2183 (
            .O(N__20844),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__2182 (
            .O(N__20841),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2181 (
            .O(N__20838),
            .I(N__20835));
    LocalMux I__2180 (
            .O(N__20835),
            .I(N__20832));
    Span4Mux_h I__2179 (
            .O(N__20832),
            .I(N__20829));
    Odrv4 I__2178 (
            .O(N__20829),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__2177 (
            .O(N__20826),
            .I(N__20823));
    InMux I__2176 (
            .O(N__20823),
            .I(N__20820));
    LocalMux I__2175 (
            .O(N__20820),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ));
    CascadeMux I__2174 (
            .O(N__20817),
            .I(N__20814));
    InMux I__2173 (
            .O(N__20814),
            .I(N__20811));
    LocalMux I__2172 (
            .O(N__20811),
            .I(N__20808));
    Odrv12 I__2171 (
            .O(N__20808),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    CascadeMux I__2170 (
            .O(N__20805),
            .I(N__20802));
    InMux I__2169 (
            .O(N__20802),
            .I(N__20799));
    LocalMux I__2168 (
            .O(N__20799),
            .I(N__20796));
    Odrv4 I__2167 (
            .O(N__20796),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__2166 (
            .O(N__20793),
            .I(N__20790));
    LocalMux I__2165 (
            .O(N__20790),
            .I(N__20787));
    Odrv4 I__2164 (
            .O(N__20787),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__2163 (
            .O(N__20784),
            .I(N__20781));
    LocalMux I__2162 (
            .O(N__20781),
            .I(N__20778));
    Span4Mux_h I__2161 (
            .O(N__20778),
            .I(N__20775));
    Odrv4 I__2160 (
            .O(N__20775),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__2159 (
            .O(N__20772),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__2158 (
            .O(N__20769),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__2157 (
            .O(N__20766),
            .I(bfn_2_26_0_));
    InMux I__2156 (
            .O(N__20763),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__2155 (
            .O(N__20760),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__2154 (
            .O(N__20757),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__2153 (
            .O(N__20754),
            .I(N__20751));
    LocalMux I__2152 (
            .O(N__20751),
            .I(N__20748));
    Odrv4 I__2151 (
            .O(N__20748),
            .I(N_88_i_i));
    InMux I__2150 (
            .O(N__20745),
            .I(N__20742));
    LocalMux I__2149 (
            .O(N__20742),
            .I(N__20739));
    Odrv4 I__2148 (
            .O(N__20739),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__2147 (
            .O(N__20736),
            .I(N__20733));
    LocalMux I__2146 (
            .O(N__20733),
            .I(N__20730));
    Span4Mux_v I__2145 (
            .O(N__20730),
            .I(N__20727));
    Odrv4 I__2144 (
            .O(N__20727),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__2143 (
            .O(N__20724),
            .I(N__20721));
    LocalMux I__2142 (
            .O(N__20721),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__2141 (
            .O(N__20718),
            .I(N__20715));
    LocalMux I__2140 (
            .O(N__20715),
            .I(N__20712));
    Span4Mux_h I__2139 (
            .O(N__20712),
            .I(N__20709));
    Odrv4 I__2138 (
            .O(N__20709),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__2137 (
            .O(N__20706),
            .I(N__20703));
    LocalMux I__2136 (
            .O(N__20703),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__2135 (
            .O(N__20700),
            .I(N__20697));
    LocalMux I__2134 (
            .O(N__20697),
            .I(N__20694));
    Span4Mux_h I__2133 (
            .O(N__20694),
            .I(N__20691));
    Odrv4 I__2132 (
            .O(N__20691),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__2131 (
            .O(N__20688),
            .I(N__20685));
    LocalMux I__2130 (
            .O(N__20685),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__2129 (
            .O(N__20682),
            .I(N__20679));
    LocalMux I__2128 (
            .O(N__20679),
            .I(N__20676));
    Span4Mux_h I__2127 (
            .O(N__20676),
            .I(N__20673));
    Odrv4 I__2126 (
            .O(N__20673),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__2125 (
            .O(N__20670),
            .I(N__20667));
    LocalMux I__2124 (
            .O(N__20667),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__2123 (
            .O(N__20664),
            .I(N__20661));
    LocalMux I__2122 (
            .O(N__20661),
            .I(N__20658));
    Span4Mux_h I__2121 (
            .O(N__20658),
            .I(N__20655));
    Odrv4 I__2120 (
            .O(N__20655),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__2119 (
            .O(N__20652),
            .I(N__20649));
    LocalMux I__2118 (
            .O(N__20649),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__2117 (
            .O(N__20646),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    InMux I__2116 (
            .O(N__20643),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__2115 (
            .O(N__20640),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__2114 (
            .O(N__20637),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__2113 (
            .O(N__20634),
            .I(N__20629));
    InMux I__2112 (
            .O(N__20633),
            .I(N__20626));
    InMux I__2111 (
            .O(N__20632),
            .I(N__20623));
    LocalMux I__2110 (
            .O(N__20629),
            .I(N__20620));
    LocalMux I__2109 (
            .O(N__20626),
            .I(pwm_duty_input_9));
    LocalMux I__2108 (
            .O(N__20623),
            .I(pwm_duty_input_9));
    Odrv4 I__2107 (
            .O(N__20620),
            .I(pwm_duty_input_9));
    InMux I__2106 (
            .O(N__20613),
            .I(N__20609));
    InMux I__2105 (
            .O(N__20612),
            .I(N__20605));
    LocalMux I__2104 (
            .O(N__20609),
            .I(N__20602));
    InMux I__2103 (
            .O(N__20608),
            .I(N__20599));
    LocalMux I__2102 (
            .O(N__20605),
            .I(N__20594));
    Span4Mux_v I__2101 (
            .O(N__20602),
            .I(N__20594));
    LocalMux I__2100 (
            .O(N__20599),
            .I(pwm_duty_input_6));
    Odrv4 I__2099 (
            .O(N__20594),
            .I(pwm_duty_input_6));
    CascadeMux I__2098 (
            .O(N__20589),
            .I(N__20585));
    InMux I__2097 (
            .O(N__20588),
            .I(N__20581));
    InMux I__2096 (
            .O(N__20585),
            .I(N__20578));
    InMux I__2095 (
            .O(N__20584),
            .I(N__20575));
    LocalMux I__2094 (
            .O(N__20581),
            .I(N__20572));
    LocalMux I__2093 (
            .O(N__20578),
            .I(pwm_duty_input_7));
    LocalMux I__2092 (
            .O(N__20575),
            .I(pwm_duty_input_7));
    Odrv4 I__2091 (
            .O(N__20572),
            .I(pwm_duty_input_7));
    InMux I__2090 (
            .O(N__20565),
            .I(N__20562));
    LocalMux I__2089 (
            .O(N__20562),
            .I(N__20557));
    InMux I__2088 (
            .O(N__20561),
            .I(N__20552));
    InMux I__2087 (
            .O(N__20560),
            .I(N__20552));
    Span4Mux_s1_h I__2086 (
            .O(N__20557),
            .I(N__20549));
    LocalMux I__2085 (
            .O(N__20552),
            .I(pwm_duty_input_8));
    Odrv4 I__2084 (
            .O(N__20549),
            .I(pwm_duty_input_8));
    InMux I__2083 (
            .O(N__20544),
            .I(N__20539));
    InMux I__2082 (
            .O(N__20543),
            .I(N__20534));
    InMux I__2081 (
            .O(N__20542),
            .I(N__20534));
    LocalMux I__2080 (
            .O(N__20539),
            .I(N__20531));
    LocalMux I__2079 (
            .O(N__20534),
            .I(pwm_duty_input_3));
    Odrv4 I__2078 (
            .O(N__20531),
            .I(pwm_duty_input_3));
    InMux I__2077 (
            .O(N__20526),
            .I(N__20521));
    InMux I__2076 (
            .O(N__20525),
            .I(N__20516));
    InMux I__2075 (
            .O(N__20524),
            .I(N__20516));
    LocalMux I__2074 (
            .O(N__20521),
            .I(N__20513));
    LocalMux I__2073 (
            .O(N__20516),
            .I(pwm_duty_input_4));
    Odrv4 I__2072 (
            .O(N__20513),
            .I(pwm_duty_input_4));
    CascadeMux I__2071 (
            .O(N__20508),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ));
    CascadeMux I__2070 (
            .O(N__20505),
            .I(N__20501));
    InMux I__2069 (
            .O(N__20504),
            .I(N__20498));
    InMux I__2068 (
            .O(N__20501),
            .I(N__20494));
    LocalMux I__2067 (
            .O(N__20498),
            .I(N__20491));
    InMux I__2066 (
            .O(N__20497),
            .I(N__20488));
    LocalMux I__2065 (
            .O(N__20494),
            .I(N__20483));
    Span4Mux_v I__2064 (
            .O(N__20491),
            .I(N__20483));
    LocalMux I__2063 (
            .O(N__20488),
            .I(pwm_duty_input_5));
    Odrv4 I__2062 (
            .O(N__20483),
            .I(pwm_duty_input_5));
    InMux I__2061 (
            .O(N__20478),
            .I(N__20475));
    LocalMux I__2060 (
            .O(N__20475),
            .I(N__20472));
    Span4Mux_h I__2059 (
            .O(N__20472),
            .I(N__20469));
    Odrv4 I__2058 (
            .O(N__20469),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__2057 (
            .O(N__20466),
            .I(N__20463));
    LocalMux I__2056 (
            .O(N__20463),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__2055 (
            .O(N__20460),
            .I(N__20457));
    LocalMux I__2054 (
            .O(N__20457),
            .I(N__20454));
    Span4Mux_v I__2053 (
            .O(N__20454),
            .I(N__20451));
    Odrv4 I__2052 (
            .O(N__20451),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__2051 (
            .O(N__20448),
            .I(N__20445));
    LocalMux I__2050 (
            .O(N__20445),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__2049 (
            .O(N__20442),
            .I(N__20439));
    LocalMux I__2048 (
            .O(N__20439),
            .I(N__20436));
    Span4Mux_h I__2047 (
            .O(N__20436),
            .I(N__20433));
    Odrv4 I__2046 (
            .O(N__20433),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__2045 (
            .O(N__20430),
            .I(N__20427));
    LocalMux I__2044 (
            .O(N__20427),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__2043 (
            .O(N__20424),
            .I(N__20421));
    LocalMux I__2042 (
            .O(N__20421),
            .I(N__20418));
    Span4Mux_h I__2041 (
            .O(N__20418),
            .I(N__20415));
    Odrv4 I__2040 (
            .O(N__20415),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__2039 (
            .O(N__20412),
            .I(N__20409));
    LocalMux I__2038 (
            .O(N__20409),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__2037 (
            .O(N__20406),
            .I(N__20403));
    LocalMux I__2036 (
            .O(N__20403),
            .I(N__20400));
    Span4Mux_v I__2035 (
            .O(N__20400),
            .I(N__20397));
    Odrv4 I__2034 (
            .O(N__20397),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__2033 (
            .O(N__20394),
            .I(N__20391));
    LocalMux I__2032 (
            .O(N__20391),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    CascadeMux I__2031 (
            .O(N__20388),
            .I(\current_shift_inst.PI_CTRL.N_31_cascade_ ));
    InMux I__2030 (
            .O(N__20385),
            .I(N__20382));
    LocalMux I__2029 (
            .O(N__20382),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__2028 (
            .O(N__20379),
            .I(\current_shift_inst.PI_CTRL.N_98_cascade_ ));
    InMux I__2027 (
            .O(N__20376),
            .I(N__20357));
    InMux I__2026 (
            .O(N__20375),
            .I(N__20357));
    InMux I__2025 (
            .O(N__20374),
            .I(N__20357));
    InMux I__2024 (
            .O(N__20373),
            .I(N__20357));
    InMux I__2023 (
            .O(N__20372),
            .I(N__20357));
    InMux I__2022 (
            .O(N__20371),
            .I(N__20357));
    InMux I__2021 (
            .O(N__20370),
            .I(N__20354));
    LocalMux I__2020 (
            .O(N__20357),
            .I(N__20351));
    LocalMux I__2019 (
            .O(N__20354),
            .I(N__20348));
    Odrv4 I__2018 (
            .O(N__20351),
            .I(\current_shift_inst.PI_CTRL.N_158 ));
    Odrv4 I__2017 (
            .O(N__20348),
            .I(\current_shift_inst.PI_CTRL.N_158 ));
    InMux I__2016 (
            .O(N__20343),
            .I(N__20340));
    LocalMux I__2015 (
            .O(N__20340),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    CascadeMux I__2014 (
            .O(N__20337),
            .I(\current_shift_inst.PI_CTRL.N_96_cascade_ ));
    InMux I__2013 (
            .O(N__20334),
            .I(N__20325));
    InMux I__2012 (
            .O(N__20333),
            .I(N__20325));
    InMux I__2011 (
            .O(N__20332),
            .I(N__20325));
    LocalMux I__2010 (
            .O(N__20325),
            .I(\current_shift_inst.PI_CTRL.N_160 ));
    InMux I__2009 (
            .O(N__20322),
            .I(N__20318));
    InMux I__2008 (
            .O(N__20321),
            .I(N__20315));
    LocalMux I__2007 (
            .O(N__20318),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    LocalMux I__2006 (
            .O(N__20315),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    InMux I__2005 (
            .O(N__20310),
            .I(N__20304));
    InMux I__2004 (
            .O(N__20309),
            .I(N__20304));
    LocalMux I__2003 (
            .O(N__20304),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__2002 (
            .O(N__20301),
            .I(N__20296));
    InMux I__2001 (
            .O(N__20300),
            .I(N__20289));
    InMux I__2000 (
            .O(N__20299),
            .I(N__20289));
    InMux I__1999 (
            .O(N__20296),
            .I(N__20282));
    InMux I__1998 (
            .O(N__20295),
            .I(N__20282));
    InMux I__1997 (
            .O(N__20294),
            .I(N__20282));
    LocalMux I__1996 (
            .O(N__20289),
            .I(N__20275));
    LocalMux I__1995 (
            .O(N__20282),
            .I(N__20275));
    InMux I__1994 (
            .O(N__20281),
            .I(N__20269));
    InMux I__1993 (
            .O(N__20280),
            .I(N__20269));
    Span4Mux_v I__1992 (
            .O(N__20275),
            .I(N__20266));
    InMux I__1991 (
            .O(N__20274),
            .I(N__20263));
    LocalMux I__1990 (
            .O(N__20269),
            .I(N__20260));
    Odrv4 I__1989 (
            .O(N__20266),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    LocalMux I__1988 (
            .O(N__20263),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    Odrv4 I__1987 (
            .O(N__20260),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    InMux I__1986 (
            .O(N__20253),
            .I(N__20250));
    LocalMux I__1985 (
            .O(N__20250),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__1984 (
            .O(N__20247),
            .I(N__20243));
    InMux I__1983 (
            .O(N__20246),
            .I(N__20240));
    LocalMux I__1982 (
            .O(N__20243),
            .I(N__20237));
    LocalMux I__1981 (
            .O(N__20240),
            .I(pwm_duty_input_1));
    Odrv4 I__1980 (
            .O(N__20237),
            .I(pwm_duty_input_1));
    InMux I__1979 (
            .O(N__20232),
            .I(N__20228));
    CascadeMux I__1978 (
            .O(N__20231),
            .I(N__20225));
    LocalMux I__1977 (
            .O(N__20228),
            .I(N__20222));
    InMux I__1976 (
            .O(N__20225),
            .I(N__20219));
    Span4Mux_v I__1975 (
            .O(N__20222),
            .I(N__20216));
    LocalMux I__1974 (
            .O(N__20219),
            .I(pwm_duty_input_2));
    Odrv4 I__1973 (
            .O(N__20216),
            .I(pwm_duty_input_2));
    InMux I__1972 (
            .O(N__20211),
            .I(N__20207));
    InMux I__1971 (
            .O(N__20210),
            .I(N__20204));
    LocalMux I__1970 (
            .O(N__20207),
            .I(N__20201));
    LocalMux I__1969 (
            .O(N__20204),
            .I(pwm_duty_input_0));
    Odrv4 I__1968 (
            .O(N__20201),
            .I(pwm_duty_input_0));
    InMux I__1967 (
            .O(N__20196),
            .I(N__20193));
    LocalMux I__1966 (
            .O(N__20193),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_1Z0Z_0 ));
    CascadeMux I__1965 (
            .O(N__20190),
            .I(\pwm_generator_inst.N_7_cascade_ ));
    CascadeMux I__1964 (
            .O(N__20187),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__1963 (
            .O(N__20184),
            .I(N__20181));
    LocalMux I__1962 (
            .O(N__20181),
            .I(N__20178));
    Odrv4 I__1961 (
            .O(N__20178),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ));
    InMux I__1960 (
            .O(N__20175),
            .I(N__20172));
    LocalMux I__1959 (
            .O(N__20172),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__1958 (
            .O(N__20169),
            .I(N__20166));
    LocalMux I__1957 (
            .O(N__20166),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__1956 (
            .O(N__20163),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ));
    InMux I__1955 (
            .O(N__20160),
            .I(N__20157));
    LocalMux I__1954 (
            .O(N__20157),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__1953 (
            .O(N__20154),
            .I(N__20151));
    LocalMux I__1952 (
            .O(N__20151),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__1951 (
            .O(N__20148),
            .I(N__20145));
    LocalMux I__1950 (
            .O(N__20145),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__1949 (
            .O(N__20142),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    CascadeMux I__1948 (
            .O(N__20139),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ));
    InMux I__1947 (
            .O(N__20136),
            .I(N__20133));
    LocalMux I__1946 (
            .O(N__20133),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    InMux I__1945 (
            .O(N__20130),
            .I(N__20127));
    LocalMux I__1944 (
            .O(N__20127),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__1943 (
            .O(N__20124),
            .I(N__20121));
    LocalMux I__1942 (
            .O(N__20121),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__1941 (
            .O(N__20118),
            .I(N__20115));
    LocalMux I__1940 (
            .O(N__20115),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    CascadeMux I__1939 (
            .O(N__20112),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ));
    InMux I__1938 (
            .O(N__20109),
            .I(N__20106));
    LocalMux I__1937 (
            .O(N__20106),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    InMux I__1936 (
            .O(N__20103),
            .I(N__20100));
    LocalMux I__1935 (
            .O(N__20100),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__1934 (
            .O(N__20097),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ));
    InMux I__1933 (
            .O(N__20094),
            .I(N__20091));
    LocalMux I__1932 (
            .O(N__20091),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    InMux I__1931 (
            .O(N__20088),
            .I(N__20085));
    LocalMux I__1930 (
            .O(N__20085),
            .I(\current_shift_inst.PI_CTRL.N_77 ));
    CascadeMux I__1929 (
            .O(N__20082),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ));
    InMux I__1928 (
            .O(N__20079),
            .I(N__20076));
    LocalMux I__1927 (
            .O(N__20076),
            .I(N__20073));
    Odrv4 I__1926 (
            .O(N__20073),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__1925 (
            .O(N__20070),
            .I(N__20067));
    LocalMux I__1924 (
            .O(N__20067),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    CascadeMux I__1923 (
            .O(N__20064),
            .I(\current_shift_inst.PI_CTRL.N_43_cascade_ ));
    InMux I__1922 (
            .O(N__20061),
            .I(N__20058));
    LocalMux I__1921 (
            .O(N__20058),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ));
    CascadeMux I__1920 (
            .O(N__20055),
            .I(N__20052));
    InMux I__1919 (
            .O(N__20052),
            .I(N__20049));
    LocalMux I__1918 (
            .O(N__20049),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__1917 (
            .O(N__20046),
            .I(N__20043));
    InMux I__1916 (
            .O(N__20043),
            .I(N__20040));
    LocalMux I__1915 (
            .O(N__20040),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__1914 (
            .O(N__20037),
            .I(N__20034));
    LocalMux I__1913 (
            .O(N__20034),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__1912 (
            .O(N__20031),
            .I(N__20028));
    LocalMux I__1911 (
            .O(N__20028),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    CascadeMux I__1910 (
            .O(N__20025),
            .I(N__20022));
    InMux I__1909 (
            .O(N__20022),
            .I(N__20019));
    LocalMux I__1908 (
            .O(N__20019),
            .I(N__20016));
    Odrv4 I__1907 (
            .O(N__20016),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__1906 (
            .O(N__20013),
            .I(N__20010));
    LocalMux I__1905 (
            .O(N__20010),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    CascadeMux I__1904 (
            .O(N__20007),
            .I(N__20004));
    InMux I__1903 (
            .O(N__20004),
            .I(N__20001));
    LocalMux I__1902 (
            .O(N__20001),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__1901 (
            .O(N__19998),
            .I(N__19995));
    LocalMux I__1900 (
            .O(N__19995),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__1899 (
            .O(N__19992),
            .I(N__19989));
    LocalMux I__1898 (
            .O(N__19989),
            .I(un7_start_stop));
    InMux I__1897 (
            .O(N__19986),
            .I(N__19983));
    LocalMux I__1896 (
            .O(N__19983),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__1895 (
            .O(N__19980),
            .I(N__19976));
    CascadeMux I__1894 (
            .O(N__19979),
            .I(N__19973));
    InMux I__1893 (
            .O(N__19976),
            .I(N__19970));
    InMux I__1892 (
            .O(N__19973),
            .I(N__19967));
    LocalMux I__1891 (
            .O(N__19970),
            .I(N__19962));
    LocalMux I__1890 (
            .O(N__19967),
            .I(N__19962));
    Span4Mux_v I__1889 (
            .O(N__19962),
            .I(N__19959));
    Span4Mux_v I__1888 (
            .O(N__19959),
            .I(N__19956));
    Odrv4 I__1887 (
            .O(N__19956),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    InMux I__1886 (
            .O(N__19953),
            .I(N__19950));
    LocalMux I__1885 (
            .O(N__19950),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__1884 (
            .O(N__19947),
            .I(N__19944));
    LocalMux I__1883 (
            .O(N__19944),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__1882 (
            .O(N__19941),
            .I(N__19938));
    LocalMux I__1881 (
            .O(N__19938),
            .I(N__19935));
    Odrv4 I__1880 (
            .O(N__19935),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__1879 (
            .O(N__19932),
            .I(N__19929));
    LocalMux I__1878 (
            .O(N__19929),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__1877 (
            .O(N__19926),
            .I(N__19923));
    LocalMux I__1876 (
            .O(N__19923),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__1875 (
            .O(N__19920),
            .I(N__19917));
    LocalMux I__1874 (
            .O(N__19917),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__1873 (
            .O(N__19914),
            .I(N__19911));
    LocalMux I__1872 (
            .O(N__19911),
            .I(N__19908));
    Odrv12 I__1871 (
            .O(N__19908),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    CascadeMux I__1870 (
            .O(N__19905),
            .I(N__19902));
    InMux I__1869 (
            .O(N__19902),
            .I(N__19899));
    LocalMux I__1868 (
            .O(N__19899),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__1867 (
            .O(N__19896),
            .I(N__19893));
    LocalMux I__1866 (
            .O(N__19893),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__1865 (
            .O(N__19890),
            .I(N__19887));
    InMux I__1864 (
            .O(N__19887),
            .I(N__19884));
    LocalMux I__1863 (
            .O(N__19884),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    CascadeMux I__1862 (
            .O(N__19881),
            .I(N__19878));
    InMux I__1861 (
            .O(N__19878),
            .I(N__19875));
    LocalMux I__1860 (
            .O(N__19875),
            .I(N__19872));
    Odrv12 I__1859 (
            .O(N__19872),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__1858 (
            .O(N__19869),
            .I(N__19866));
    LocalMux I__1857 (
            .O(N__19866),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    CascadeMux I__1856 (
            .O(N__19863),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ));
    CascadeMux I__1855 (
            .O(N__19860),
            .I(N__19857));
    InMux I__1854 (
            .O(N__19857),
            .I(N__19854));
    LocalMux I__1853 (
            .O(N__19854),
            .I(N__19851));
    Odrv12 I__1852 (
            .O(N__19851),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__1851 (
            .O(N__19848),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__1850 (
            .O(N__19845),
            .I(N__19842));
    InMux I__1849 (
            .O(N__19842),
            .I(N__19839));
    LocalMux I__1848 (
            .O(N__19839),
            .I(N__19836));
    Span4Mux_v I__1847 (
            .O(N__19836),
            .I(N__19833));
    Odrv4 I__1846 (
            .O(N__19833),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__1845 (
            .O(N__19830),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__1844 (
            .O(N__19827),
            .I(N__19824));
    InMux I__1843 (
            .O(N__19824),
            .I(N__19821));
    LocalMux I__1842 (
            .O(N__19821),
            .I(N__19818));
    Span4Mux_v I__1841 (
            .O(N__19818),
            .I(N__19815));
    Odrv4 I__1840 (
            .O(N__19815),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__1839 (
            .O(N__19812),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__1838 (
            .O(N__19809),
            .I(N__19806));
    InMux I__1837 (
            .O(N__19806),
            .I(N__19803));
    LocalMux I__1836 (
            .O(N__19803),
            .I(N__19800));
    Span4Mux_v I__1835 (
            .O(N__19800),
            .I(N__19797));
    Odrv4 I__1834 (
            .O(N__19797),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__1833 (
            .O(N__19794),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__1832 (
            .O(N__19791),
            .I(N__19788));
    InMux I__1831 (
            .O(N__19788),
            .I(N__19785));
    LocalMux I__1830 (
            .O(N__19785),
            .I(N__19782));
    Span4Mux_v I__1829 (
            .O(N__19782),
            .I(N__19779));
    Odrv4 I__1828 (
            .O(N__19779),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__1827 (
            .O(N__19776),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__1826 (
            .O(N__19773),
            .I(N__19770));
    LocalMux I__1825 (
            .O(N__19770),
            .I(N__19767));
    Odrv12 I__1824 (
            .O(N__19767),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    CascadeMux I__1823 (
            .O(N__19764),
            .I(N__19761));
    InMux I__1822 (
            .O(N__19761),
            .I(N__19758));
    LocalMux I__1821 (
            .O(N__19758),
            .I(N__19755));
    Odrv12 I__1820 (
            .O(N__19755),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    InMux I__1819 (
            .O(N__19752),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__1818 (
            .O(N__19749),
            .I(N__19746));
    LocalMux I__1817 (
            .O(N__19746),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    CascadeMux I__1816 (
            .O(N__19743),
            .I(N__19740));
    InMux I__1815 (
            .O(N__19740),
            .I(N__19737));
    LocalMux I__1814 (
            .O(N__19737),
            .I(N__19734));
    Odrv4 I__1813 (
            .O(N__19734),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__1812 (
            .O(N__19731),
            .I(bfn_1_14_0_));
    CascadeMux I__1811 (
            .O(N__19728),
            .I(N__19725));
    InMux I__1810 (
            .O(N__19725),
            .I(N__19722));
    LocalMux I__1809 (
            .O(N__19722),
            .I(N__19719));
    Span4Mux_v I__1808 (
            .O(N__19719),
            .I(N__19716));
    Odrv4 I__1807 (
            .O(N__19716),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__1806 (
            .O(N__19713),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__1805 (
            .O(N__19710),
            .I(N__19707));
    InMux I__1804 (
            .O(N__19707),
            .I(N__19704));
    LocalMux I__1803 (
            .O(N__19704),
            .I(N__19701));
    Span4Mux_v I__1802 (
            .O(N__19701),
            .I(N__19698));
    Odrv4 I__1801 (
            .O(N__19698),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__1800 (
            .O(N__19695),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__1799 (
            .O(N__19692),
            .I(N__19689));
    LocalMux I__1798 (
            .O(N__19689),
            .I(N__19686));
    Span4Mux_v I__1797 (
            .O(N__19686),
            .I(N__19683));
    Odrv4 I__1796 (
            .O(N__19683),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__1795 (
            .O(N__19680),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__1794 (
            .O(N__19677),
            .I(N__19674));
    InMux I__1793 (
            .O(N__19674),
            .I(N__19671));
    LocalMux I__1792 (
            .O(N__19671),
            .I(N__19668));
    Span4Mux_v I__1791 (
            .O(N__19668),
            .I(N__19665));
    Odrv4 I__1790 (
            .O(N__19665),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__1789 (
            .O(N__19662),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__1788 (
            .O(N__19659),
            .I(N__19656));
    InMux I__1787 (
            .O(N__19656),
            .I(N__19653));
    LocalMux I__1786 (
            .O(N__19653),
            .I(N__19650));
    Span4Mux_v I__1785 (
            .O(N__19650),
            .I(N__19647));
    Odrv4 I__1784 (
            .O(N__19647),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__1783 (
            .O(N__19644),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    InMux I__1782 (
            .O(N__19641),
            .I(N__19638));
    LocalMux I__1781 (
            .O(N__19638),
            .I(N__19635));
    Odrv12 I__1780 (
            .O(N__19635),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__1779 (
            .O(N__19632),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__1778 (
            .O(N__19629),
            .I(N__19626));
    InMux I__1777 (
            .O(N__19626),
            .I(N__19623));
    LocalMux I__1776 (
            .O(N__19623),
            .I(N__19620));
    Odrv12 I__1775 (
            .O(N__19620),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__1774 (
            .O(N__19617),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    InMux I__1773 (
            .O(N__19614),
            .I(N__19611));
    LocalMux I__1772 (
            .O(N__19611),
            .I(N__19608));
    Span4Mux_v I__1771 (
            .O(N__19608),
            .I(N__19605));
    Odrv4 I__1770 (
            .O(N__19605),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__1769 (
            .O(N__19602),
            .I(bfn_1_15_0_));
    CascadeMux I__1768 (
            .O(N__19599),
            .I(N__19596));
    InMux I__1767 (
            .O(N__19596),
            .I(N__19593));
    LocalMux I__1766 (
            .O(N__19593),
            .I(N__19590));
    Span4Mux_v I__1765 (
            .O(N__19590),
            .I(N__19587));
    Span4Mux_v I__1764 (
            .O(N__19587),
            .I(N__19584));
    Odrv4 I__1763 (
            .O(N__19584),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__1762 (
            .O(N__19581),
            .I(bfn_1_13_0_));
    CascadeMux I__1761 (
            .O(N__19578),
            .I(N__19575));
    InMux I__1760 (
            .O(N__19575),
            .I(N__19572));
    LocalMux I__1759 (
            .O(N__19572),
            .I(N__19569));
    Span4Mux_v I__1758 (
            .O(N__19569),
            .I(N__19566));
    Span4Mux_v I__1757 (
            .O(N__19566),
            .I(N__19563));
    Odrv4 I__1756 (
            .O(N__19563),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__1755 (
            .O(N__19560),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__1754 (
            .O(N__19557),
            .I(N__19554));
    InMux I__1753 (
            .O(N__19554),
            .I(N__19551));
    LocalMux I__1752 (
            .O(N__19551),
            .I(N__19548));
    Span4Mux_v I__1751 (
            .O(N__19548),
            .I(N__19545));
    Odrv4 I__1750 (
            .O(N__19545),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__1749 (
            .O(N__19542),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    CascadeMux I__1748 (
            .O(N__19539),
            .I(N__19536));
    InMux I__1747 (
            .O(N__19536),
            .I(N__19533));
    LocalMux I__1746 (
            .O(N__19533),
            .I(N__19530));
    Span4Mux_v I__1745 (
            .O(N__19530),
            .I(N__19527));
    Odrv4 I__1744 (
            .O(N__19527),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__1743 (
            .O(N__19524),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__1742 (
            .O(N__19521),
            .I(N__19518));
    InMux I__1741 (
            .O(N__19518),
            .I(N__19515));
    LocalMux I__1740 (
            .O(N__19515),
            .I(N__19512));
    Span4Mux_v I__1739 (
            .O(N__19512),
            .I(N__19509));
    Odrv4 I__1738 (
            .O(N__19509),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__1737 (
            .O(N__19506),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    CascadeMux I__1736 (
            .O(N__19503),
            .I(N__19500));
    InMux I__1735 (
            .O(N__19500),
            .I(N__19497));
    LocalMux I__1734 (
            .O(N__19497),
            .I(N__19494));
    Span4Mux_v I__1733 (
            .O(N__19494),
            .I(N__19491));
    Odrv4 I__1732 (
            .O(N__19491),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__1731 (
            .O(N__19488),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__1730 (
            .O(N__19485),
            .I(N__19482));
    InMux I__1729 (
            .O(N__19482),
            .I(N__19479));
    LocalMux I__1728 (
            .O(N__19479),
            .I(N__19476));
    Span4Mux_v I__1727 (
            .O(N__19476),
            .I(N__19473));
    Odrv4 I__1726 (
            .O(N__19473),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__1725 (
            .O(N__19470),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__1724 (
            .O(N__19467),
            .I(N__19464));
    InMux I__1723 (
            .O(N__19464),
            .I(N__19461));
    LocalMux I__1722 (
            .O(N__19461),
            .I(N__19458));
    Odrv12 I__1721 (
            .O(N__19458),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__1720 (
            .O(N__19455),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    CascadeMux I__1719 (
            .O(N__19452),
            .I(N__19449));
    InMux I__1718 (
            .O(N__19449),
            .I(N__19446));
    LocalMux I__1717 (
            .O(N__19446),
            .I(N__19443));
    Span4Mux_v I__1716 (
            .O(N__19443),
            .I(N__19440));
    Odrv4 I__1715 (
            .O(N__19440),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    CascadeMux I__1714 (
            .O(N__19437),
            .I(N__19434));
    InMux I__1713 (
            .O(N__19434),
            .I(N__19431));
    LocalMux I__1712 (
            .O(N__19431),
            .I(N__19428));
    Span4Mux_v I__1711 (
            .O(N__19428),
            .I(N__19425));
    Span4Mux_v I__1710 (
            .O(N__19425),
            .I(N__19422));
    Odrv4 I__1709 (
            .O(N__19422),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__1708 (
            .O(N__19419),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    CascadeMux I__1707 (
            .O(N__19416),
            .I(N__19413));
    InMux I__1706 (
            .O(N__19413),
            .I(N__19410));
    LocalMux I__1705 (
            .O(N__19410),
            .I(N__19407));
    Span4Mux_v I__1704 (
            .O(N__19407),
            .I(N__19404));
    Odrv4 I__1703 (
            .O(N__19404),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__1702 (
            .O(N__19401),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    InMux I__1701 (
            .O(N__19398),
            .I(N__19395));
    LocalMux I__1700 (
            .O(N__19395),
            .I(N__19392));
    Span4Mux_v I__1699 (
            .O(N__19392),
            .I(N__19389));
    Odrv4 I__1698 (
            .O(N__19389),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    InMux I__1697 (
            .O(N__19386),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    InMux I__1696 (
            .O(N__19383),
            .I(N__19380));
    LocalMux I__1695 (
            .O(N__19380),
            .I(N__19377));
    Span4Mux_v I__1694 (
            .O(N__19377),
            .I(N__19374));
    Odrv4 I__1693 (
            .O(N__19374),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__1692 (
            .O(N__19371),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__1691 (
            .O(N__19368),
            .I(N__19365));
    InMux I__1690 (
            .O(N__19365),
            .I(N__19362));
    LocalMux I__1689 (
            .O(N__19362),
            .I(N__19359));
    Span4Mux_v I__1688 (
            .O(N__19359),
            .I(N__19356));
    Odrv4 I__1687 (
            .O(N__19356),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__1686 (
            .O(N__19353),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__1685 (
            .O(N__19350),
            .I(N__19347));
    InMux I__1684 (
            .O(N__19347),
            .I(N__19344));
    LocalMux I__1683 (
            .O(N__19344),
            .I(N__19341));
    Span4Mux_v I__1682 (
            .O(N__19341),
            .I(N__19338));
    Odrv4 I__1681 (
            .O(N__19338),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__1680 (
            .O(N__19335),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__1679 (
            .O(N__19332),
            .I(N__19329));
    InMux I__1678 (
            .O(N__19329),
            .I(N__19326));
    LocalMux I__1677 (
            .O(N__19326),
            .I(N__19323));
    Span4Mux_v I__1676 (
            .O(N__19323),
            .I(N__19320));
    Odrv4 I__1675 (
            .O(N__19320),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__1674 (
            .O(N__19317),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    InMux I__1673 (
            .O(N__19314),
            .I(N__19311));
    LocalMux I__1672 (
            .O(N__19311),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__1671 (
            .O(N__19308),
            .I(bfn_1_10_0_));
    InMux I__1670 (
            .O(N__19305),
            .I(N__19302));
    LocalMux I__1669 (
            .O(N__19302),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__1668 (
            .O(N__19299),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__1667 (
            .O(N__19296),
            .I(N__19293));
    LocalMux I__1666 (
            .O(N__19293),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__1665 (
            .O(N__19290),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__1664 (
            .O(N__19287),
            .I(N__19284));
    LocalMux I__1663 (
            .O(N__19284),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__1662 (
            .O(N__19281),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__1661 (
            .O(N__19278),
            .I(N__19275));
    LocalMux I__1660 (
            .O(N__19275),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__1659 (
            .O(N__19272),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__1658 (
            .O(N__19269),
            .I(N__19266));
    LocalMux I__1657 (
            .O(N__19266),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__1656 (
            .O(N__19263),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__1655 (
            .O(N__19260),
            .I(N__19257));
    LocalMux I__1654 (
            .O(N__19257),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    InMux I__1653 (
            .O(N__19254),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__1652 (
            .O(N__19251),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    InMux I__1651 (
            .O(N__19248),
            .I(N__19245));
    LocalMux I__1650 (
            .O(N__19245),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__1649 (
            .O(N__19242),
            .I(N__19228));
    CascadeMux I__1648 (
            .O(N__19241),
            .I(N__19225));
    CascadeMux I__1647 (
            .O(N__19240),
            .I(N__19222));
    CascadeMux I__1646 (
            .O(N__19239),
            .I(N__19219));
    CascadeMux I__1645 (
            .O(N__19238),
            .I(N__19216));
    CascadeMux I__1644 (
            .O(N__19237),
            .I(N__19213));
    CascadeMux I__1643 (
            .O(N__19236),
            .I(N__19210));
    CascadeMux I__1642 (
            .O(N__19235),
            .I(N__19207));
    CascadeMux I__1641 (
            .O(N__19234),
            .I(N__19204));
    CascadeMux I__1640 (
            .O(N__19233),
            .I(N__19201));
    CascadeMux I__1639 (
            .O(N__19232),
            .I(N__19198));
    CascadeMux I__1638 (
            .O(N__19231),
            .I(N__19195));
    LocalMux I__1637 (
            .O(N__19228),
            .I(N__19192));
    InMux I__1636 (
            .O(N__19225),
            .I(N__19185));
    InMux I__1635 (
            .O(N__19222),
            .I(N__19185));
    InMux I__1634 (
            .O(N__19219),
            .I(N__19185));
    InMux I__1633 (
            .O(N__19216),
            .I(N__19176));
    InMux I__1632 (
            .O(N__19213),
            .I(N__19176));
    InMux I__1631 (
            .O(N__19210),
            .I(N__19176));
    InMux I__1630 (
            .O(N__19207),
            .I(N__19176));
    InMux I__1629 (
            .O(N__19204),
            .I(N__19171));
    InMux I__1628 (
            .O(N__19201),
            .I(N__19171));
    InMux I__1627 (
            .O(N__19198),
            .I(N__19166));
    InMux I__1626 (
            .O(N__19195),
            .I(N__19166));
    Span4Mux_v I__1625 (
            .O(N__19192),
            .I(N__19155));
    LocalMux I__1624 (
            .O(N__19185),
            .I(N__19155));
    LocalMux I__1623 (
            .O(N__19176),
            .I(N__19155));
    LocalMux I__1622 (
            .O(N__19171),
            .I(N__19155));
    LocalMux I__1621 (
            .O(N__19166),
            .I(N__19155));
    Odrv4 I__1620 (
            .O(N__19155),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    InMux I__1619 (
            .O(N__19152),
            .I(N__19149));
    LocalMux I__1618 (
            .O(N__19149),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__1617 (
            .O(N__19146),
            .I(N__19143));
    InMux I__1616 (
            .O(N__19143),
            .I(N__19140));
    LocalMux I__1615 (
            .O(N__19140),
            .I(N__19137));
    Odrv4 I__1614 (
            .O(N__19137),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    InMux I__1613 (
            .O(N__19134),
            .I(N__19131));
    LocalMux I__1612 (
            .O(N__19131),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__1611 (
            .O(N__19128),
            .I(N__19125));
    InMux I__1610 (
            .O(N__19125),
            .I(N__19122));
    LocalMux I__1609 (
            .O(N__19122),
            .I(N__19119));
    Odrv4 I__1608 (
            .O(N__19119),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    InMux I__1607 (
            .O(N__19116),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__1606 (
            .O(N__19113),
            .I(N__19110));
    LocalMux I__1605 (
            .O(N__19110),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__1604 (
            .O(N__19107),
            .I(N__19104));
    InMux I__1603 (
            .O(N__19104),
            .I(N__19101));
    LocalMux I__1602 (
            .O(N__19101),
            .I(N__19098));
    Odrv4 I__1601 (
            .O(N__19098),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    InMux I__1600 (
            .O(N__19095),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    InMux I__1599 (
            .O(N__19092),
            .I(N__19089));
    LocalMux I__1598 (
            .O(N__19089),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__1597 (
            .O(N__19086),
            .I(N__19083));
    InMux I__1596 (
            .O(N__19083),
            .I(N__19080));
    LocalMux I__1595 (
            .O(N__19080),
            .I(N__19077));
    Odrv4 I__1594 (
            .O(N__19077),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__1593 (
            .O(N__19074),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    InMux I__1592 (
            .O(N__19071),
            .I(N__19068));
    LocalMux I__1591 (
            .O(N__19068),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__1590 (
            .O(N__19065),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    InMux I__1589 (
            .O(N__19062),
            .I(N__19059));
    LocalMux I__1588 (
            .O(N__19059),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__1587 (
            .O(N__19056),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__1586 (
            .O(N__19053),
            .I(N__19050));
    LocalMux I__1585 (
            .O(N__19050),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__1584 (
            .O(N__19047),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    InMux I__1583 (
            .O(N__19044),
            .I(N__19041));
    LocalMux I__1582 (
            .O(N__19041),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__1581 (
            .O(N__19038),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    IoInMux I__1580 (
            .O(N__19035),
            .I(N__19032));
    LocalMux I__1579 (
            .O(N__19032),
            .I(N__19029));
    Span4Mux_s3_v I__1578 (
            .O(N__19029),
            .I(N__19026));
    Span4Mux_h I__1577 (
            .O(N__19026),
            .I(N__19023));
    Sp12to4 I__1576 (
            .O(N__19023),
            .I(N__19020));
    Span12Mux_v I__1575 (
            .O(N__19020),
            .I(N__19017));
    Span12Mux_v I__1574 (
            .O(N__19017),
            .I(N__19014));
    Odrv12 I__1573 (
            .O(N__19014),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1572 (
            .O(N__19011),
            .I(N__19008));
    LocalMux I__1571 (
            .O(N__19008),
            .I(N__19005));
    IoSpan4Mux I__1570 (
            .O(N__19005),
            .I(N__19002));
    IoSpan4Mux I__1569 (
            .O(N__19002),
            .I(N__18999));
    Odrv4 I__1568 (
            .O(N__18999),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_4_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_22_0_));
    defparam IN_MUX_bfv_4_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_23_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_4_23_0_));
    defparam IN_MUX_bfv_4_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_24_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_4_24_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_5_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_23_0_));
    defparam IN_MUX_bfv_5_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_24_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_5_24_0_));
    defparam IN_MUX_bfv_5_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_25_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_5_25_0_));
    defparam IN_MUX_bfv_3_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_24_0_));
    defparam IN_MUX_bfv_3_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_25_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_3_25_0_));
    defparam IN_MUX_bfv_2_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_24_0_));
    defparam IN_MUX_bfv_2_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_25_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_2_25_0_));
    defparam IN_MUX_bfv_2_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_26_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_2_26_0_));
    defparam IN_MUX_bfv_8_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_24_0_));
    defparam IN_MUX_bfv_8_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_25_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_8_25_0_));
    defparam IN_MUX_bfv_7_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_26_0_));
    defparam IN_MUX_bfv_7_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_27_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_7_27_0_));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_15 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_23 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_17_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_25_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_17_25_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_9_16_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19035),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19011),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__34794),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_161_i_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__33684),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__41286),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__38678),
            .CLKHFEN(N__38680),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__38679),
            .RGB2PWM(N__20754),
            .RGB1(rgb_g),
            .CURREN(N__38848),
            .RGB2(rgb_b),
            .RGB1PWM(N__19992),
            .RGB0PWM(N__49479),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__19152),
            .in2(N__19146),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__19134),
            .in2(N__19128),
            .in3(N__19116),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__19113),
            .in2(N__19107),
            .in3(N__19095),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__19092),
            .in2(N__19086),
            .in3(N__19074),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__19071),
            .in2(N__19231),
            .in3(N__19065),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__19062),
            .in2(N__19233),
            .in3(N__19056),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(N__19053),
            .in2(N__19232),
            .in3(N__19047),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(N__19044),
            .in2(N__19234),
            .in3(N__19038),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__19314),
            .in2(N__19235),
            .in3(N__19308),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__19305),
            .in2(N__19239),
            .in3(N__19299),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__19296),
            .in2(N__19236),
            .in3(N__19290),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__19287),
            .in2(N__19240),
            .in3(N__19281),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__19278),
            .in2(N__19237),
            .in3(N__19272),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__19269),
            .in2(N__19241),
            .in3(N__19263),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__19260),
            .in2(N__19238),
            .in3(N__19254),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19251),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__19248),
            .in2(_gnd_net_),
            .in3(N__19242),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__21113),
            .in2(N__19979),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__21067),
            .in2(N__19437),
            .in3(N__19419),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__21012),
            .in2(N__19416),
            .in3(N__19401),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__19398),
            .in2(N__20930),
            .in3(N__19386),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__19383),
            .in2(N__22670),
            .in3(N__19371),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__21509),
            .in2(N__19368),
            .in3(N__19353),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__21453),
            .in2(N__19350),
            .in3(N__19335),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(N__21430),
            .in2(N__19332),
            .in3(N__19317),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__21376),
            .in2(N__19599),
            .in3(N__19581),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__22917),
            .in2(N__19578),
            .in3(N__19560),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__21307),
            .in2(N__19557),
            .in3(N__19542),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__21253),
            .in2(N__19539),
            .in3(N__19524),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__22965),
            .in2(N__19521),
            .in3(N__19506),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__21858),
            .in2(N__19503),
            .in3(N__19488),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__23007),
            .in2(N__19485),
            .in3(N__19470),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__22882),
            .in2(N__19467),
            .in3(N__19455),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__21774),
            .in2(N__19452),
            .in3(N__19731),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__21718),
            .in2(N__19728),
            .in3(N__19713),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__21663),
            .in2(N__19710),
            .in3(N__19695),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__19692),
            .in2(N__21619),
            .in3(N__19680),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__21558),
            .in2(N__19677),
            .in3(N__19662),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__22302),
            .in2(N__19659),
            .in3(N__19644),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__19641),
            .in2(N__22247),
            .in3(N__19632),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__22182),
            .in2(N__19629),
            .in3(N__19617),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__19614),
            .in2(N__22136),
            .in3(N__19602),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__22075),
            .in2(N__19860),
            .in3(N__19848),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__22017),
            .in2(N__19845),
            .in3(N__19830),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__21963),
            .in2(N__19827),
            .in3(N__19812),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__21908),
            .in2(N__19809),
            .in3(N__19794),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__22590),
            .in2(N__19791),
            .in3(N__19776),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6  (
            .in0(N__19773),
            .in1(N__23506),
            .in2(N__19764),
            .in3(N__19752),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_2 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_2  (
            .in0(N__23519),
            .in1(N__23203),
            .in2(N__23378),
            .in3(N__19749),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49901),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_16_3 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_1_16_3  (
            .in0(N__23201),
            .in1(N__23522),
            .in2(N__19743),
            .in3(N__23339),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49901),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5  (
            .in0(N__23202),
            .in1(N__23523),
            .in2(N__19905),
            .in3(N__23340),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49901),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_6 .LUT_INIT=16'b1111111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_6  (
            .in0(N__23520),
            .in1(N__23204),
            .in2(N__23379),
            .in3(N__19896),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49901),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_7 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_7  (
            .in0(N__23200),
            .in1(N__23521),
            .in2(N__19890),
            .in3(N__23338),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49901),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_1_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_1_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_1_17_2 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_1_17_2  (
            .in0(N__23524),
            .in1(N__23369),
            .in2(N__19881),
            .in3(N__23230),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49888),
            .ce(),
            .sr(N__49441));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_1_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_1_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_1_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28734),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49878),
            .ce(),
            .sr(N__49444));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__21155),
            .in2(_gnd_net_),
            .in3(N__21137),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49878),
            .ce(),
            .sr(N__49444));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_1_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_1_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__21807),
            .in2(_gnd_net_),
            .in3(N__21828),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_1_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_1_20_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_1_20_5  (
            .in0(N__22104),
            .in1(N__19869),
            .in2(N__22275),
            .in3(N__22050),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_1_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_1_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_1_20_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_1_20_6  (
            .in0(N__20118),
            .in1(N__20148),
            .in2(N__19863),
            .in3(N__20103),
            .lcout(\current_shift_inst.PI_CTRL.N_158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_0 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_0  (
            .in0(N__29782),
            .in1(N__20371),
            .in2(N__22386),
            .in3(N__20299),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_22_1 .LUT_INIT=16'b1010000011111100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_22_1  (
            .in0(N__20372),
            .in1(N__20294),
            .in2(N__22515),
            .in3(N__29783),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2  (
            .in0(N__29784),
            .in1(N__20373),
            .in2(N__22422),
            .in3(N__20300),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_3 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_3  (
            .in0(N__20979),
            .in1(N__20343),
            .in2(_gnd_net_),
            .in3(N__20322),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_4 .LUT_INIT=16'b1101110101010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_4  (
            .in0(N__29786),
            .in1(N__20375),
            .in2(N__20301),
            .in3(N__22484),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_22_5 .LUT_INIT=16'b1011001110110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_22_5  (
            .in0(N__20374),
            .in1(N__29785),
            .in2(N__22455),
            .in3(N__20295),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_7 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_7  (
            .in0(N__20376),
            .in1(N__20895),
            .in2(N__22347),
            .in3(N__20385),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(N__49453));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(N__21039),
            .in2(_gnd_net_),
            .in3(N__20334),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49825),
            .ce(),
            .sr(N__49454));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_23_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_23_3  (
            .in0(N__20333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19914),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49825),
            .ce(),
            .sr(N__49454));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(N__22527),
            .in2(_gnd_net_),
            .in3(N__20332),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49825),
            .ce(),
            .sr(N__49454));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_24_1  (
            .in0(N__23897),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23915),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un7_start_stop_LC_1_29_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.un7_start_stop_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un7_start_stop_LC_1_29_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.un7_start_stop_LC_1_29_0  (
            .in0(N__49478),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35106),
            .lcout(un7_start_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_2_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_2_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_2_12_2 .LUT_INIT=16'b1111001100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_2_12_2  (
            .in0(N__23388),
            .in1(N__23578),
            .in2(N__23241),
            .in3(N__19986),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49935),
            .ce(),
            .sr(N__49418));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_3 .LUT_INIT=16'b0101101001001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_3  (
            .in0(N__21123),
            .in1(N__23390),
            .in2(N__19980),
            .in3(N__23213),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49935),
            .ce(),
            .sr(N__49418));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_2_12_7 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_2_12_7  (
            .in0(N__19953),
            .in1(N__23389),
            .in2(_gnd_net_),
            .in3(N__23212),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49935),
            .ce(),
            .sr(N__49418));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_2_13_3 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_2_13_3  (
            .in0(N__23387),
            .in1(N__23586),
            .in2(N__23243),
            .in3(N__19947),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49924),
            .ce(),
            .sr(N__49422));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_0 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_0  (
            .in0(N__23423),
            .in1(N__23585),
            .in2(N__23239),
            .in3(N__19941),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49427));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1  (
            .in0(N__23581),
            .in1(N__23426),
            .in2(N__23245),
            .in3(N__19932),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49427));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_2_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_2_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_2_14_2 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_2_14_2  (
            .in0(N__23420),
            .in1(N__23582),
            .in2(N__23237),
            .in3(N__19926),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49427));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_3 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_3  (
            .in0(N__23580),
            .in1(N__23425),
            .in2(N__23244),
            .in3(N__19920),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49427));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_4 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_4  (
            .in0(N__23422),
            .in1(N__23584),
            .in2(N__20055),
            .in3(N__23223),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49427));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_5 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_5  (
            .in0(N__23579),
            .in1(N__23424),
            .in2(N__20046),
            .in3(N__23196),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49427));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_6 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_6  (
            .in0(N__23421),
            .in1(N__23583),
            .in2(N__23238),
            .in3(N__20037),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(),
            .sr(N__49427));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1 .LUT_INIT=16'b1100111111001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1  (
            .in0(N__23371),
            .in1(N__20031),
            .in2(N__23207),
            .in3(N__23529),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_2_15_4 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_2_15_4  (
            .in0(N__23525),
            .in1(N__23373),
            .in2(N__20025),
            .in3(N__23150),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5  (
            .in0(N__23370),
            .in1(N__23527),
            .in2(N__23206),
            .in3(N__20013),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_6 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_6  (
            .in0(N__23526),
            .in1(N__23374),
            .in2(N__20007),
            .in3(N__23149),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_7 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_7  (
            .in0(N__23372),
            .in1(N__23528),
            .in2(N__23208),
            .in3(N__19998),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_16_0  (
            .in0(N__21906),
            .in1(N__23008),
            .in2(N__22938),
            .in3(N__22973),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_16_3  (
            .in0(N__21670),
            .in1(N__21717),
            .in2(N__22316),
            .in3(N__21779),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_16_4  (
            .in0(N__21907),
            .in1(N__22240),
            .in2(N__20097),
            .in3(N__20094),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_16_5 .LUT_INIT=16'b0000000101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_16_5  (
            .in0(N__20929),
            .in1(N__21136),
            .in2(N__21075),
            .in3(N__21017),
            .lcout(\current_shift_inst.PI_CTRL.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_16_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_16_6  (
            .in0(N__21016),
            .in1(N__20928),
            .in2(N__20826),
            .in3(N__22668),
            .lcout(\current_shift_inst.PI_CTRL.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_2  (
            .in0(N__22883),
            .in1(N__21868),
            .in2(N__21249),
            .in3(N__21311),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_17_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__22068),
            .in2(_gnd_net_),
            .in3(N__21559),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5  (
            .in0(N__21432),
            .in1(N__22669),
            .in2(_gnd_net_),
            .in3(N__21469),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_6 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_6  (
            .in0(N__21508),
            .in1(N__20088),
            .in2(N__20082),
            .in3(N__21380),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_7  (
            .in0(N__20079),
            .in1(N__20070),
            .in2(N__20064),
            .in3(N__20136),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_0  (
            .in0(N__21618),
            .in1(N__20130),
            .in2(N__22190),
            .in3(N__20061),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_1  (
            .in0(N__20124),
            .in1(N__23530),
            .in2(N__20139),
            .in3(N__22239),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_3  (
            .in0(N__22594),
            .in1(N__22018),
            .in2(N__21974),
            .in3(N__22135),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_5  (
            .in0(N__21719),
            .in1(N__21674),
            .in2(N__22315),
            .in3(N__21778),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_0  (
            .in0(N__21194),
            .in1(N__22155),
            .in2(N__22208),
            .in3(N__21839),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_19_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(N__22265),
            .in2(_gnd_net_),
            .in3(N__21530),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_2  (
            .in0(N__21329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21209),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_19_3  (
            .in0(N__21840),
            .in1(N__21639),
            .in2(N__21588),
            .in3(N__21195),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_4  (
            .in0(N__21531),
            .in1(N__21888),
            .in2(N__22209),
            .in3(N__22154),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_5  (
            .in0(N__21279),
            .in1(N__21936),
            .in2(N__20112),
            .in3(N__20109),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6  (
            .in0(N__21800),
            .in1(N__21887),
            .in2(N__21330),
            .in3(N__21821),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_19_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_19_7  (
            .in0(N__21278),
            .in1(N__21210),
            .in2(N__20187),
            .in3(N__20154),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_20_2  (
            .in0(N__22100),
            .in1(N__21584),
            .in2(N__22049),
            .in3(N__21638),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_2_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_2_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_2_20_3  (
            .in0(N__20184),
            .in1(N__21935),
            .in2(N__22562),
            .in3(N__21989),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_4  (
            .in0(N__20175),
            .in1(N__20169),
            .in2(N__20163),
            .in3(N__20160),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_5  (
            .in0(_gnd_net_),
            .in1(N__21749),
            .in2(_gnd_net_),
            .in3(N__21692),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_7  (
            .in0(N__21693),
            .in1(N__21750),
            .in2(N__22563),
            .in3(N__21990),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_3  (
            .in0(_gnd_net_),
            .in1(N__22480),
            .in2(_gnd_net_),
            .in3(N__22375),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_4  (
            .in0(N__22448),
            .in1(N__22511),
            .in2(N__20142),
            .in3(N__22415),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(\current_shift_inst.PI_CTRL.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_21_5 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_21_5  (
            .in0(N__29758),
            .in1(N__20890),
            .in2(N__20388),
            .in3(N__20274),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_22_0  (
            .in0(_gnd_net_),
            .in1(N__20889),
            .in2(_gnd_net_),
            .in3(N__20974),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_1 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_1  (
            .in0(N__29764),
            .in1(N__22340),
            .in2(N__20379),
            .in3(N__20370),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(\current_shift_inst.PI_CTRL.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_22_2 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_22_2  (
            .in0(N__20975),
            .in1(N__20253),
            .in2(N__20337),
            .in3(N__20321),
            .lcout(\current_shift_inst.PI_CTRL.N_160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_22_5 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_22_5  (
            .in0(N__29763),
            .in1(N__20309),
            .in2(N__20894),
            .in3(N__20281),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_1_0_LC_2_22_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_1_0_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_1_0_LC_2_22_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_1_0_LC_2_22_6  (
            .in0(N__20612),
            .in1(N__20584),
            .in2(N__20505),
            .in3(N__20632),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_7  (
            .in0(N__29762),
            .in1(N__20310),
            .in2(_gnd_net_),
            .in3(N__20280),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o2_1_LC_2_23_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o2_1_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o2_1_LC_2_23_1 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o2_1_LC_2_23_1  (
            .in0(N__20246),
            .in1(N__20543),
            .in2(N__20231),
            .in3(N__20210),
            .lcout(),
            .ltout(\pwm_generator_inst.N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_2 .LUT_INIT=16'b1101110111111101;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_2  (
            .in0(N__20561),
            .in1(N__20196),
            .in2(N__20190),
            .in3(N__20524),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3  (
            .in0(N__20633),
            .in1(N__20608),
            .in2(N__20589),
            .in3(N__20560),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_23_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_23_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_23_4  (
            .in0(N__20542),
            .in1(N__20525),
            .in2(N__20508),
            .in3(N__20497),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(N__20466),
            .in2(_gnd_net_),
            .in3(N__20478),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_2_24_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_24_1  (
            .in0(_gnd_net_),
            .in1(N__20448),
            .in2(_gnd_net_),
            .in3(N__20460),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_24_2  (
            .in0(_gnd_net_),
            .in1(N__20430),
            .in2(_gnd_net_),
            .in3(N__20442),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_24_3  (
            .in0(_gnd_net_),
            .in1(N__20412),
            .in2(_gnd_net_),
            .in3(N__20424),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_24_4  (
            .in0(_gnd_net_),
            .in1(N__20394),
            .in2(_gnd_net_),
            .in3(N__20406),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(N__20724),
            .in2(_gnd_net_),
            .in3(N__20736),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(N__20706),
            .in2(_gnd_net_),
            .in3(N__20718),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_24_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_24_7  (
            .in0(_gnd_net_),
            .in1(N__20688),
            .in2(_gnd_net_),
            .in3(N__20700),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_25_0  (
            .in0(_gnd_net_),
            .in1(N__20670),
            .in2(_gnd_net_),
            .in3(N__20682),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_2_25_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_25_1  (
            .in0(_gnd_net_),
            .in1(N__20652),
            .in2(_gnd_net_),
            .in3(N__20664),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_25_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_25_2  (
            .in0(_gnd_net_),
            .in1(N__23893),
            .in2(_gnd_net_),
            .in3(N__20646),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_25_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_25_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_25_3  (
            .in0(N__24745),
            .in1(N__23841),
            .in2(_gnd_net_),
            .in3(N__20643),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_25_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_25_4  (
            .in0(_gnd_net_),
            .in1(N__23966),
            .in2(_gnd_net_),
            .in3(N__20640),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_25_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_25_5  (
            .in0(_gnd_net_),
            .in1(N__24093),
            .in2(_gnd_net_),
            .in3(N__20637),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_25_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_25_6  (
            .in0(_gnd_net_),
            .in1(N__24122),
            .in2(_gnd_net_),
            .in3(N__20772),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_25_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_25_7  (
            .in0(_gnd_net_),
            .in1(N__22784),
            .in2(_gnd_net_),
            .in3(N__20769),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_26_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_26_0  (
            .in0(_gnd_net_),
            .in1(N__22810),
            .in2(_gnd_net_),
            .in3(N__20766),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_26_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_26_1  (
            .in0(_gnd_net_),
            .in1(N__22719),
            .in2(_gnd_net_),
            .in3(N__20763),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_26_2  (
            .in0(_gnd_net_),
            .in1(N__22757),
            .in2(_gnd_net_),
            .in3(N__20760),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_26_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20757),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_7  (
            .in0(N__22758),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23715),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.N_88_i_i_LC_2_30_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_88_i_i_LC_2_30_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_88_i_i_LC_2_30_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \phase_controller_inst1.N_88_i_i_LC_2_30_1  (
            .in0(N__35105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49477),
            .lcout(N_88_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_1  (
            .in0(N__20745),
            .in1(N__23418),
            .in2(_gnd_net_),
            .in3(N__23221),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49925),
            .ce(),
            .sr(N__49414));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_3 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_3  (
            .in0(N__23598),
            .in1(N__23419),
            .in2(N__20817),
            .in3(N__23222),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49925),
            .ce(),
            .sr(N__49414));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29213),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49913),
            .ce(),
            .sr(N__49419));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_13_3 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_3_13_3  (
            .in0(N__23592),
            .in1(N__23381),
            .in2(N__20805),
            .in3(N__23217),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49913),
            .ce(),
            .sr(N__49419));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(N__29192),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49913),
            .ce(),
            .sr(N__49419));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_13_6 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_3_13_6  (
            .in0(N__23380),
            .in1(N__23593),
            .in2(N__23242),
            .in3(N__20793),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49913),
            .ce(),
            .sr(N__49419));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_3_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_3_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_3_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_3_13_7  (
            .in0(N__28688),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49913),
            .ce(),
            .sr(N__49419));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_1 .LUT_INIT=16'b1010000010101011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_1  (
            .in0(N__20784),
            .in1(N__23427),
            .in2(N__23240),
            .in3(N__23597),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49423));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28664),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49423));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29102),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49423));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_3_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_3_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_3_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30803),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49903),
            .ce(),
            .sr(N__49423));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29327),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49428));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29244),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49428));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_3_15_3 .LUT_INIT=16'b1100110001000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_3_15_3  (
            .in0(N__23591),
            .in1(N__20838),
            .in2(N__23417),
            .in3(N__23151),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49428));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_4  (
            .in0(N__29678),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49428));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29072),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49428));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_3_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_3_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_3_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29009),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49890),
            .ce(),
            .sr(N__49428));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_1  (
            .in0(N__21423),
            .in1(N__21495),
            .in2(N__21470),
            .in3(N__21366),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_2  (
            .in0(N__23552),
            .in1(N__22186),
            .in2(N__21566),
            .in3(N__21620),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_3  (
            .in0(N__22076),
            .in1(N__22019),
            .in2(N__21970),
            .in3(N__22128),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(N__21872),
            .in2(_gnd_net_),
            .in3(N__21306),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_5  (
            .in0(N__22595),
            .in1(N__21257),
            .in2(N__21183),
            .in3(N__22848),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_6  (
            .in0(N__21180),
            .in1(N__21174),
            .in2(N__21168),
            .in3(N__21165),
            .lcout(\current_shift_inst.PI_CTRL.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__21159),
            .in2(N__21141),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__21087),
            .in2(N__21074),
            .in3(N__21024),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49435));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__21021),
            .in2(N__20991),
            .in3(N__20946),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49435));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__20943),
            .in2(N__20934),
            .in3(N__20856),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49435));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__20853),
            .in2(N__22671),
            .in3(N__20841),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49435));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__21519),
            .in2(N__21510),
            .in3(N__21474),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49435));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__23619),
            .in2(N__21471),
            .in3(N__21435),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49435));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__23049),
            .in2(N__21431),
            .in3(N__21396),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__49866),
            .ce(),
            .sr(N__49435));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__21393),
            .in2(N__21384),
            .in3(N__21342),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49439));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__21339),
            .in2(N__22934),
            .in3(N__21318),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49439));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(N__22842),
            .in2(N__21315),
            .in3(N__21270),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49439));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__21267),
            .in2(N__21258),
            .in3(N__21198),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49439));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__23040),
            .in2(N__22977),
            .in3(N__21186),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49439));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__22836),
            .in2(N__21876),
            .in3(N__21831),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49439));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__23028),
            .in2(N__23016),
            .in3(N__21810),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49439));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__23679),
            .in2(N__22890),
            .in3(N__21789),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49439));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__24045),
            .in2(N__21786),
            .in3(N__21741),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__49843),
            .ce(),
            .sr(N__49442));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__21738),
            .in2(N__21726),
            .in3(N__21681),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__49843),
            .ce(),
            .sr(N__49442));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__23640),
            .in2(N__21678),
            .in3(N__21627),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__49843),
            .ce(),
            .sr(N__49442));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__21624),
            .in2(N__23634),
            .in3(N__21573),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__49843),
            .ce(),
            .sr(N__49442));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__22542),
            .in2(N__21570),
            .in3(N__21522),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__49843),
            .ce(),
            .sr(N__49442));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__22329),
            .in2(N__22320),
            .in3(N__22254),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__49843),
            .ce(),
            .sr(N__49442));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__23652),
            .in2(N__22251),
            .in3(N__22194),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__49843),
            .ce(),
            .sr(N__49442));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__22191),
            .in2(N__23691),
            .in3(N__22146),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__49843),
            .ce(),
            .sr(N__49442));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__23673),
            .in2(N__22143),
            .in3(N__22089),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__49833),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__23625),
            .in2(N__22086),
            .in3(N__22032),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__49833),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__23646),
            .in2(N__22029),
            .in3(N__21981),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__49833),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__24033),
            .in2(N__21978),
            .in3(N__21924),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__49833),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__23664),
            .in2(N__21921),
            .in3(N__21879),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__49833),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(N__24018),
            .in2(N__22602),
            .in3(N__22548),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__49833),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6  (
            .in0(N__23590),
            .in1(N__29796),
            .in2(_gnd_net_),
            .in3(N__22545),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49833),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_3_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_3_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_3_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_3_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29712),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49833),
            .ce(),
            .sr(N__49445));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22536),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49826),
            .ce(),
            .sr(N__49450));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_22_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_22_2  (
            .in0(_gnd_net_),
            .in1(N__22504),
            .in2(_gnd_net_),
            .in3(N__22485),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_3  (
            .in0(N__22447),
            .in1(N__22414),
            .in2(N__22389),
            .in3(N__22382),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_3_23_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_3_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_3_23_1  (
            .in0(_gnd_net_),
            .in1(N__22717),
            .in2(_gnd_net_),
            .in3(N__23729),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_3_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_3_23_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_3_23_3  (
            .in0(_gnd_net_),
            .in1(N__23765),
            .in2(_gnd_net_),
            .in3(N__22783),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_3_23_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_3_23_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_3_23_4  (
            .in0(_gnd_net_),
            .in1(N__23939),
            .in2(_gnd_net_),
            .in3(N__23965),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_23_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_23_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_23_5  (
            .in0(N__24146),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24121),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_24_0  (
            .in0(_gnd_net_),
            .in1(N__23865),
            .in2(N__24771),
            .in3(N__24770),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ),
            .ltout(),
            .carryin(bfn_3_24_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_24_1  (
            .in0(_gnd_net_),
            .in1(N__22629),
            .in2(_gnd_net_),
            .in3(N__22623),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_24_2  (
            .in0(_gnd_net_),
            .in1(N__23928),
            .in2(_gnd_net_),
            .in3(N__22620),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_24_3  (
            .in0(_gnd_net_),
            .in1(N__24051),
            .in2(_gnd_net_),
            .in3(N__22617),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_24_4  (
            .in0(_gnd_net_),
            .in1(N__24099),
            .in2(_gnd_net_),
            .in3(N__22614),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_24_5  (
            .in0(_gnd_net_),
            .in1(N__22764),
            .in2(_gnd_net_),
            .in3(N__22611),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_24_6  (
            .in0(_gnd_net_),
            .in1(N__22797),
            .in2(_gnd_net_),
            .in3(N__22608),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_24_7  (
            .in0(_gnd_net_),
            .in1(N__22692),
            .in2(_gnd_net_),
            .in3(N__22605),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_25_0  (
            .in0(_gnd_net_),
            .in1(N__22731),
            .in2(_gnd_net_),
            .in3(N__22830),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ),
            .ltout(),
            .carryin(bfn_3_25_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_25_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_25_1  (
            .in0(N__24755),
            .in1(N__22827),
            .in2(N__23859),
            .in3(N__22821),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_3_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_3_25_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_3_25_2  (
            .in0(N__22812),
            .in1(_gnd_net_),
            .in2(N__23751),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_25_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_25_3 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_25_3  (
            .in0(N__22818),
            .in1(N__23750),
            .in2(N__24765),
            .in3(N__22811),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_25_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_25_5 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_25_5  (
            .in0(N__22791),
            .in1(N__22785),
            .in2(N__24764),
            .in3(N__23772),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_3_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_3_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_3_25_6 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_3_25_6  (
            .in0(N__24757),
            .in1(N__22756),
            .in2(N__22743),
            .in3(N__23714),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_3_25_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_3_25_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_3_25_7  (
            .in0(N__23733),
            .in1(N__22725),
            .in2(N__24766),
            .in3(N__22718),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_13_1 .LUT_INIT=16'b1010001010100011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_4_13_1  (
            .in0(N__22686),
            .in1(N__23588),
            .in2(N__23247),
            .in3(N__23430),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(),
            .sr(N__49415));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29162),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(),
            .sr(N__49415));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_4_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_4_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_4_13_7 .LUT_INIT=16'b1010111110101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_4_13_7  (
            .in0(N__23607),
            .in1(N__23429),
            .in2(N__23246),
            .in3(N__23589),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(),
            .sr(N__49415));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_4_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_4_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_4_14_0 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_4_14_0  (
            .in0(N__23587),
            .in1(N__23428),
            .in2(N__23262),
            .in3(N__23205),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49891),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29135),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49891),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29468),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49891),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_4_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_4_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_4_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29411),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49891),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_16_6  (
            .in0(N__23012),
            .in1(N__22969),
            .in2(N__22933),
            .in3(N__22881),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29039),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29444),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_4_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29628),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_4_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_4_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_4_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29390),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49844),
            .ce(),
            .sr(N__49436));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_4_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_4_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_4_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_4_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29594),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49844),
            .ce(),
            .sr(N__49436));
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_4_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_4_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_29_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29865),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49844),
            .ce(),
            .sr(N__49436));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_4_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_4_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_4_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29655),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(N__49440));
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_4_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_4_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_4_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_27_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29531),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(N__49440));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_4_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_4_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_4_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29303),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(N__49440));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_4_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29271),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(N__49440));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_4_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_4_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_4_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_4_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29564),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49827),
            .ce(),
            .sr(N__49443));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_4_22_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_4_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_4_22_0  (
            .in0(_gnd_net_),
            .in1(N__23840),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_22_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_4_22_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_4_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_4_22_1  (
            .in0(_gnd_net_),
            .in1(N__23817),
            .in2(_gnd_net_),
            .in3(N__23805),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_4_22_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_4_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_4_22_2  (
            .in0(_gnd_net_),
            .in1(N__23802),
            .in2(_gnd_net_),
            .in3(N__23790),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_4_22_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_4_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_4_22_3  (
            .in0(_gnd_net_),
            .in1(N__23787),
            .in2(_gnd_net_),
            .in3(N__23775),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_4_22_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_4_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_4_22_4  (
            .in0(_gnd_net_),
            .in1(N__24399),
            .in2(_gnd_net_),
            .in3(N__23754),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_4_22_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_4_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_4_22_5  (
            .in0(_gnd_net_),
            .in1(N__24357),
            .in2(N__38572),
            .in3(N__23736),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_4_22_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_4_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_4_22_6  (
            .in0(_gnd_net_),
            .in1(N__38531),
            .in2(N__24315),
            .in3(N__23718),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_4_22_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_4_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_4_22_7  (
            .in0(_gnd_net_),
            .in1(N__24273),
            .in2(N__38573),
            .in3(N__23694),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_4_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_4_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_4_23_0  (
            .in0(_gnd_net_),
            .in1(N__24237),
            .in2(_gnd_net_),
            .in3(N__23844),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_4_23_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_4_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_4_23_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_4_23_1  (
            .in0(_gnd_net_),
            .in1(N__24198),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_4_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_4_23_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_4_23_2  (
            .in0(_gnd_net_),
            .in1(N__24159),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_4_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_4_23_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_4_23_3  (
            .in0(_gnd_net_),
            .in1(N__24660),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_4_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_4_23_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_4_23_4  (
            .in0(_gnd_net_),
            .in1(N__24615),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_4_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_4_23_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_4_23_5  (
            .in0(_gnd_net_),
            .in1(N__24570),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_4_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_4_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_4_23_6  (
            .in0(_gnd_net_),
            .in1(N__24540),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_4_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_4_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_4_23_7  (
            .in0(_gnd_net_),
            .in1(N__24516),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_4_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_4_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_4_24_0  (
            .in0(_gnd_net_),
            .in1(N__24492),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_24_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_4_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_4_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__24471),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_4_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_4_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_4_24_2  (
            .in0(_gnd_net_),
            .in1(N__24441),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_4_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_4_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_4_24_3  (
            .in0(_gnd_net_),
            .in1(N__24789),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_4_24_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_4_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_4_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24006),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_24_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_24_5 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_24_5  (
            .in0(N__26984),
            .in1(N__24003),
            .in2(N__48870),
            .in3(N__26918),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_24_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_24_7 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_24_7  (
            .in0(N__26983),
            .in1(N__23997),
            .in2(N__48869),
            .in3(N__26917),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_25_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_25_0 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_25_0  (
            .in0(N__26989),
            .in1(N__48780),
            .in2(N__23991),
            .in3(N__26919),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_4_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_4_25_1 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_4_25_1  (
            .in0(N__24737),
            .in1(N__23979),
            .in2(N__23970),
            .in3(N__23943),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_2  (
            .in0(N__23922),
            .in1(N__23904),
            .in2(N__23877),
            .in3(N__24736),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_3 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_3  (
            .in0(N__24738),
            .in1(N__24150),
            .in2(N__24135),
            .in3(N__24123),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_25_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_25_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_25_5  (
            .in0(N__24092),
            .in1(_gnd_net_),
            .in2(N__24066),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_6 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_6  (
            .in0(N__24756),
            .in1(N__24078),
            .in2(N__24069),
            .in3(N__24065),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_5_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_5_6_5 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_5_6_5  (
            .in0(N__25782),
            .in1(N__28194),
            .in2(N__25763),
            .in3(N__28221),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_5_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_5_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_5_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_5_7_5  (
            .in0(N__24852),
            .in1(N__26397),
            .in2(_gnd_net_),
            .in3(N__36681),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49950),
            .ce(N__33338),
            .sr(N__49384));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29357),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49867),
            .ce(),
            .sr(N__49421));
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_28_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29492),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49857),
            .ce(),
            .sr(N__49424));
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_5_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_30_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29834),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49835),
            .ce(),
            .sr(N__49432));
    defparam CONSTANT_ONE_LUT4_LC_5_22_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_22_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_22_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_5_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_5_23_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_5_23_0  (
            .in0(_gnd_net_),
            .in1(N__24432),
            .in2(N__24417),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_5_23_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_5_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_5_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_5_23_1  (
            .in0(_gnd_net_),
            .in1(N__24393),
            .in2(N__24375),
            .in3(N__24351),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_5_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_5_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_5_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_5_23_2  (
            .in0(_gnd_net_),
            .in1(N__24348),
            .in2(N__24333),
            .in3(N__24306),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_5_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_5_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_5_23_3  (
            .in0(_gnd_net_),
            .in1(N__24303),
            .in2(N__24288),
            .in3(N__24267),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_5_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_5_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_5_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_5_23_4  (
            .in0(_gnd_net_),
            .in1(N__24264),
            .in2(N__24252),
            .in3(N__24231),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_5_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_5_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_5_23_5  (
            .in0(_gnd_net_),
            .in1(N__24228),
            .in2(N__24216),
            .in3(N__24192),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_5_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_5_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_5_23_6  (
            .in0(_gnd_net_),
            .in1(N__24189),
            .in2(N__24174),
            .in3(N__24153),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_5_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_5_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_5_23_7  (
            .in0(_gnd_net_),
            .in1(N__24690),
            .in2(N__24675),
            .in3(N__24654),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_5_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_5_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_5_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_5_24_0  (
            .in0(_gnd_net_),
            .in1(N__24651),
            .in2(N__24636),
            .in3(N__24609),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_5_24_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_5_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_5_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_5_24_1  (
            .in0(_gnd_net_),
            .in1(N__24606),
            .in2(N__24591),
            .in3(N__24564),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_5_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_5_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_5_24_2  (
            .in0(_gnd_net_),
            .in1(N__48936),
            .in2(N__24561),
            .in3(N__24534),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_5_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_5_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_5_24_3  (
            .in0(_gnd_net_),
            .in1(N__24531),
            .in2(N__48951),
            .in3(N__24510),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_5_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_5_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_5_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_5_24_4  (
            .in0(_gnd_net_),
            .in1(N__48940),
            .in2(N__24507),
            .in3(N__24486),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_5_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_5_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_5_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_5_24_5  (
            .in0(_gnd_net_),
            .in1(N__24483),
            .in2(N__48952),
            .in3(N__24465),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_5_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_5_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_5_24_6  (
            .in0(_gnd_net_),
            .in1(N__48944),
            .in2(N__24462),
            .in3(N__24435),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_5_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_5_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_5_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_5_24_7  (
            .in0(_gnd_net_),
            .in1(N__48663),
            .in2(N__48953),
            .in3(N__24783),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_5_25_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_5_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_5_25_0  (
            .in0(N__24780),
            .in1(N__30693),
            .in2(_gnd_net_),
            .in3(N__24774),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_7_2_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_7_2_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_7_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_7_2_3  (
            .in0(N__24896),
            .in1(N__25994),
            .in2(_gnd_net_),
            .in3(N__36649),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(N__31249),
            .sr(N__49340));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_7_2_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_7_2_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_7_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_7_2_4  (
            .in0(N__36645),
            .in1(N__24848),
            .in2(_gnd_net_),
            .in3(N__26396),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(N__31249),
            .sr(N__49340));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_7_2_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_7_2_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_7_2_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_7_2_6  (
            .in0(N__26142),
            .in1(_gnd_net_),
            .in2(N__36703),
            .in3(N__24913),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(N__31249),
            .sr(N__49340));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_2_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_2_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_2_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_7_2_7  (
            .in0(N__30228),
            .in1(N__30185),
            .in2(_gnd_net_),
            .in3(N__36650),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(N__31249),
            .sr(N__49340));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_7_3_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_7_3_0 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_7_3_0  (
            .in0(N__24824),
            .in1(N__28076),
            .in2(N__24809),
            .in3(N__28109),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_3_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_3_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_3_6  (
            .in0(N__24917),
            .in1(N__26141),
            .in2(_gnd_net_),
            .in3(N__36632),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_4_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_4_0  (
            .in0(N__24825),
            .in1(N__28077),
            .in2(N__24810),
            .in3(N__28110),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_7_4_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_7_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_7_4_3  (
            .in0(N__30223),
            .in1(N__30184),
            .in2(_gnd_net_),
            .in3(N__36637),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_4_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_4_6  (
            .in0(N__36636),
            .in1(N__24895),
            .in2(_gnd_net_),
            .in3(N__25998),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_7_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_7_5_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_7_5_0  (
            .in0(N__28050),
            .in1(N__25889),
            .in2(N__28029),
            .in3(N__24933),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_7_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_7_5_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_7_5_1  (
            .in0(N__24932),
            .in1(N__28024),
            .in2(N__25893),
            .in3(N__28049),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_5_5  (
            .in0(N__24847),
            .in1(N__26389),
            .in2(_gnd_net_),
            .in3(N__36651),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_7_6_1  (
            .in0(N__31307),
            .in1(N__31356),
            .in2(_gnd_net_),
            .in3(N__36602),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49946),
            .ce(N__31248),
            .sr(N__49370));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_7_6_5  (
            .in0(N__28508),
            .in1(N__28481),
            .in2(_gnd_net_),
            .in3(N__36603),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49946),
            .ce(N__31248),
            .sr(N__49370));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_7_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_7_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_7_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_7_7_2  (
            .in0(N__36545),
            .in1(N__28799),
            .in2(_gnd_net_),
            .in3(N__28776),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49936),
            .ce(N__31200),
            .sr(N__49374));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_7_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_7_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_7_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_7_7_7  (
            .in0(N__30893),
            .in1(N__30920),
            .in2(_gnd_net_),
            .in3(N__36546),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49936),
            .ce(N__31200),
            .sr(N__49374));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_7_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_7_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_7_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_7_8_2  (
            .in0(N__36469),
            .in1(N__28974),
            .in2(_gnd_net_),
            .in3(N__28936),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(N__31255),
            .sr(N__49380));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_7_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_7_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_7_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_7_8_3  (
            .in0(N__33159),
            .in1(N__33203),
            .in2(_gnd_net_),
            .in3(N__36470),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(N__31255),
            .sr(N__49380));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_7_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_7_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_7_8_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_7_8_5  (
            .in0(N__25874),
            .in1(_gnd_net_),
            .in2(N__26682),
            .in3(N__36471),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(N__31255),
            .sr(N__49380));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_7_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_7_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_7_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_7_9_1  (
            .in0(N__36464),
            .in1(N__24921),
            .in2(_gnd_net_),
            .in3(N__26140),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(N__33339),
            .sr(N__49385));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_7_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_7_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_7_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_7_9_3  (
            .in0(N__36462),
            .in1(N__26742),
            .in2(_gnd_net_),
            .in3(N__25713),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(N__33339),
            .sr(N__49385));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_7_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_7_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_7_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_7_9_4  (
            .in0(N__24897),
            .in1(N__25993),
            .in2(_gnd_net_),
            .in3(N__36465),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(N__33339),
            .sr(N__49385));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_7_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_7_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_7_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_7_9_6  (
            .in0(N__26681),
            .in1(N__25873),
            .in2(_gnd_net_),
            .in3(N__36466),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(N__33339),
            .sr(N__49385));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_7_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_7_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_7_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_7_9_7  (
            .in0(N__36463),
            .in1(N__26589),
            .in2(_gnd_net_),
            .in3(N__25635),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(N__33339),
            .sr(N__49385));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_7_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_7_10_0 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_7_10_0  (
            .in0(N__31772),
            .in1(N__24873),
            .in2(N__24864),
            .in3(N__31796),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_7_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_7_10_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_7_10_1  (
            .in0(N__24872),
            .in1(N__31773),
            .in2(N__31797),
            .in3(N__24863),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_7_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_7_11_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__25931),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49892),
            .ce(N__27061),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26240),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49892),
            .ce(N__27061),
            .sr(N__49393));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_7_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_7_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_7_11_5  (
            .in0(N__36477),
            .in1(N__28504),
            .in2(_gnd_net_),
            .in3(N__28470),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_7_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_7_12_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_7_12_2  (
            .in0(N__36478),
            .in1(N__30916),
            .in2(_gnd_net_),
            .in3(N__30889),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_13_0  (
            .in0(N__25115),
            .in1(N__25921),
            .in2(_gnd_net_),
            .in3(N__24951),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__49868),
            .ce(N__25160),
            .sr(N__49401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_13_1  (
            .in0(N__25103),
            .in1(N__26230),
            .in2(_gnd_net_),
            .in3(N__24948),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__49868),
            .ce(N__25160),
            .sr(N__49401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_13_2  (
            .in0(N__25116),
            .in1(N__26204),
            .in2(_gnd_net_),
            .in3(N__24945),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__49868),
            .ce(N__25160),
            .sr(N__49401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_13_3  (
            .in0(N__25104),
            .in1(N__26185),
            .in2(_gnd_net_),
            .in3(N__24942),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__49868),
            .ce(N__25160),
            .sr(N__49401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_13_4  (
            .in0(N__25117),
            .in1(N__26158),
            .in2(_gnd_net_),
            .in3(N__24939),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__49868),
            .ce(N__25160),
            .sr(N__49401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_13_5  (
            .in0(N__25105),
            .in1(N__26098),
            .in2(_gnd_net_),
            .in3(N__24936),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__49868),
            .ce(N__25160),
            .sr(N__49401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_13_6  (
            .in0(N__25118),
            .in1(N__26074),
            .in2(_gnd_net_),
            .in3(N__24978),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__49868),
            .ce(N__25160),
            .sr(N__49401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_13_7  (
            .in0(N__25106),
            .in1(N__26041),
            .in2(_gnd_net_),
            .in3(N__24975),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__49868),
            .ce(N__25160),
            .sr(N__49401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_14_0  (
            .in0(N__25102),
            .in1(N__26017),
            .in2(_gnd_net_),
            .in3(N__24972),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__49858),
            .ce(N__25161),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_14_1  (
            .in0(N__25114),
            .in1(N__26491),
            .in2(_gnd_net_),
            .in3(N__24969),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__49858),
            .ce(N__25161),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_14_2  (
            .in0(N__25099),
            .in1(N__26461),
            .in2(_gnd_net_),
            .in3(N__24966),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__49858),
            .ce(N__25161),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_14_3  (
            .in0(N__25111),
            .in1(N__26432),
            .in2(_gnd_net_),
            .in3(N__24963),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__49858),
            .ce(N__25161),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_14_4  (
            .in0(N__25100),
            .in1(N__26413),
            .in2(_gnd_net_),
            .in3(N__24960),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__49858),
            .ce(N__25161),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_14_5  (
            .in0(N__25112),
            .in1(N__26344),
            .in2(_gnd_net_),
            .in3(N__24957),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__49858),
            .ce(N__25161),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_14_6  (
            .in0(N__25101),
            .in1(N__26312),
            .in2(_gnd_net_),
            .in3(N__24954),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__49858),
            .ce(N__25161),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_14_7  (
            .in0(N__25113),
            .in1(N__26290),
            .in2(_gnd_net_),
            .in3(N__25005),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__49858),
            .ce(N__25161),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_15_0  (
            .in0(N__25107),
            .in1(N__26263),
            .in2(_gnd_net_),
            .in3(N__25002),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__49845),
            .ce(N__25159),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_15_1  (
            .in0(N__25119),
            .in1(N__26803),
            .in2(_gnd_net_),
            .in3(N__24999),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__49845),
            .ce(N__25159),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_15_2  (
            .in0(N__25108),
            .in1(N__26779),
            .in2(_gnd_net_),
            .in3(N__24996),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__49845),
            .ce(N__25159),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_15_3  (
            .in0(N__25120),
            .in1(N__26758),
            .in2(_gnd_net_),
            .in3(N__24993),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__49845),
            .ce(N__25159),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_15_4  (
            .in0(N__25109),
            .in1(N__26698),
            .in2(_gnd_net_),
            .in3(N__24990),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__49845),
            .ce(N__25159),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_15_5  (
            .in0(N__25121),
            .in1(N__26630),
            .in2(_gnd_net_),
            .in3(N__24987),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__49845),
            .ce(N__25159),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_15_6  (
            .in0(N__25110),
            .in1(N__26605),
            .in2(_gnd_net_),
            .in3(N__24984),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__49845),
            .ce(N__25159),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_15_7  (
            .in0(N__25122),
            .in1(N__26545),
            .in2(_gnd_net_),
            .in3(N__24981),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__49845),
            .ce(N__25159),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_16_0  (
            .in0(N__25093),
            .in1(N__26521),
            .in2(_gnd_net_),
            .in3(N__25179),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__49836),
            .ce(N__25149),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_16_1  (
            .in0(N__25097),
            .in1(N__27172),
            .in2(_gnd_net_),
            .in3(N__25176),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__49836),
            .ce(N__25149),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_16_2  (
            .in0(N__25094),
            .in1(N__27130),
            .in2(_gnd_net_),
            .in3(N__25173),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__49836),
            .ce(N__25149),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_16_3  (
            .in0(N__25098),
            .in1(N__27088),
            .in2(_gnd_net_),
            .in3(N__25170),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__49836),
            .ce(N__25149),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_16_4  (
            .in0(N__25095),
            .in1(N__27149),
            .in2(_gnd_net_),
            .in3(N__25167),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__49836),
            .ce(N__25149),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_16_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_16_5  (
            .in0(N__27107),
            .in1(N__25096),
            .in2(_gnd_net_),
            .in3(N__25164),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49836),
            .ce(N__25149),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_17_0 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_17_0  (
            .in0(N__25313),
            .in1(_gnd_net_),
            .in2(N__25296),
            .in3(N__25274),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_7_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_7_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__25312),
            .in2(_gnd_net_),
            .in3(N__25292),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_165_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25311),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_7_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_7_18_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_7_18_4  (
            .in0(N__25314),
            .in1(N__25291),
            .in2(_gnd_net_),
            .in3(N__25275),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49821),
            .ce(),
            .sr(N__49425));
    defparam \delay_measurement_inst.stop_timer_tr_LC_7_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25273),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25248),
            .ce(),
            .sr(N__49429));
    defparam \delay_measurement_inst.start_timer_tr_LC_7_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_7_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25272),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25247),
            .ce(),
            .sr(N__49433));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_7_24_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_7_24_0 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_7_24_0  (
            .in0(N__27003),
            .in1(N__25236),
            .in2(N__48852),
            .in3(N__26912),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_7_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_7_24_1 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_7_24_1  (
            .in0(N__26913),
            .in1(N__25227),
            .in2(N__48849),
            .in3(N__27004),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_7_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_7_24_2 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_7_24_2  (
            .in0(N__27002),
            .in1(N__25218),
            .in2(N__48851),
            .in3(N__26911),
            .lcout(\pwm_generator_inst.threshold_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_7_24_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_7_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_7_24_4 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_7_24_4  (
            .in0(N__27006),
            .in1(N__26915),
            .in2(N__25209),
            .in3(N__48796),
            .lcout(\pwm_generator_inst.threshold_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_7_24_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_7_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_7_24_7 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_7_24_7  (
            .in0(N__26914),
            .in1(N__27005),
            .in2(N__48850),
            .in3(N__25197),
            .lcout(\pwm_generator_inst.threshold_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_7_25_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_7_25_7 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_7_25_7  (
            .in0(N__26990),
            .in1(N__25188),
            .in2(N__48781),
            .in3(N__26916),
            .lcout(\pwm_generator_inst.threshold_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_7_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_7_26_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_7_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_7_26_0  (
            .in0(N__27402),
            .in1(N__27563),
            .in2(_gnd_net_),
            .in3(N__25341),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_26_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__49805),
            .ce(),
            .sr(N__49451));
    defparam \pwm_generator_inst.counter_1_LC_7_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_7_26_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_7_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_7_26_1  (
            .in0(N__27387),
            .in1(N__27500),
            .in2(_gnd_net_),
            .in3(N__25338),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__49805),
            .ce(),
            .sr(N__49451));
    defparam \pwm_generator_inst.counter_2_LC_7_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_7_26_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_7_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_7_26_2  (
            .in0(N__27403),
            .in1(N__27542),
            .in2(_gnd_net_),
            .in3(N__25335),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__49805),
            .ce(),
            .sr(N__49451));
    defparam \pwm_generator_inst.counter_3_LC_7_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_7_26_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_7_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_7_26_3  (
            .in0(N__27388),
            .in1(N__27476),
            .in2(_gnd_net_),
            .in3(N__25332),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__49805),
            .ce(),
            .sr(N__49451));
    defparam \pwm_generator_inst.counter_4_LC_7_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_7_26_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_7_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_7_26_4  (
            .in0(N__27404),
            .in1(N__27521),
            .in2(_gnd_net_),
            .in3(N__25329),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__49805),
            .ce(),
            .sr(N__49451));
    defparam \pwm_generator_inst.counter_5_LC_7_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_7_26_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_7_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_7_26_5  (
            .in0(N__27389),
            .in1(N__27424),
            .in2(_gnd_net_),
            .in3(N__25326),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__49805),
            .ce(),
            .sr(N__49451));
    defparam \pwm_generator_inst.counter_6_LC_7_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_7_26_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_7_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_7_26_6  (
            .in0(N__27405),
            .in1(N__27448),
            .in2(_gnd_net_),
            .in3(N__25323),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__49805),
            .ce(),
            .sr(N__49451));
    defparam \pwm_generator_inst.counter_7_LC_7_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_7_26_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_7_26_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_7_26_7  (
            .in0(N__27390),
            .in1(N__27587),
            .in2(_gnd_net_),
            .in3(N__25320),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__49805),
            .ce(),
            .sr(N__49451));
    defparam \pwm_generator_inst.counter_8_LC_7_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_7_27_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_7_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_7_27_0  (
            .in0(N__27392),
            .in1(N__27629),
            .in2(_gnd_net_),
            .in3(N__25317),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_27_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__49801),
            .ce(),
            .sr(N__49452));
    defparam \pwm_generator_inst.counter_9_LC_7_27_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_7_27_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_7_27_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_7_27_1  (
            .in0(N__27608),
            .in1(N__27391),
            .in2(_gnd_net_),
            .in3(N__25446),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49801),
            .ce(),
            .sr(N__49452));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_8_1_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_8_1_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(N__27795),
            .in2(N__25443),
            .in3(N__27778),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_8_1_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_8_1_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(N__25434),
            .in2(N__25422),
            .in3(N__27762),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_8_1_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_8_1_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__29730),
            .in2(N__25413),
            .in3(N__27744),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_8_1_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_8_1_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_8_1_3  (
            .in0(N__27726),
            .in1(N__25656),
            .in2(N__25401),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_8_1_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_8_1_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_8_1_4  (
            .in0(_gnd_net_),
            .in1(N__25392),
            .in2(N__25386),
            .in3(N__27708),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_8_1_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_8_1_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(N__27333),
            .in2(N__25374),
            .in3(N__27690),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_8_1_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_8_1_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(N__25365),
            .in2(N__25359),
            .in3(N__27672),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_8_1_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_8_1_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(N__25836),
            .in2(N__25350),
            .in3(N__27651),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_8_2_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_8_2_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__29973),
            .in2(N__25524),
            .in3(N__27930),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_8_2_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_8_2_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__25722),
            .in2(N__25515),
            .in3(N__27912),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_8_2_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_8_2_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(N__25506),
            .in2(N__25500),
            .in3(N__27894),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_8_2_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_8_2_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__25905),
            .in2(N__25491),
            .in3(N__27876),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_8_2_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_8_2_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(N__27339),
            .in2(N__25482),
            .in3(N__27858),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_8_2_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_8_2_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__31281),
            .in2(N__25470),
            .in3(N__27837),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_8_2_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_8_2_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_8_2_6  (
            .in0(N__27816),
            .in1(N__25452),
            .in2(N__25461),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_8_2_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_8_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__29961),
            .in2(N__29901),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_8_3_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_8_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__25590),
            .in2(N__25584),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_8_3_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_8_3_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__25572),
            .in2(N__25563),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_8_3_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_8_3_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__25662),
            .in2(N__25533),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_8_3_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_8_3_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__25599),
            .in2(N__25647),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_8_3_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_8_3_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__25815),
            .in2(N__25827),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_8_3_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_8_3_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(N__28173),
            .in2(N__28128),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_8_3_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_8_3_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(N__25734),
            .in2(N__25551),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_3_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25536),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_4_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_4_0  (
            .in0(N__25692),
            .in1(N__27983),
            .in2(N__25683),
            .in3(N__28001),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_8_4_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_8_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_8_4_1  (
            .in0(N__26740),
            .in1(N__36633),
            .in2(_gnd_net_),
            .in3(N__25706),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_8_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_8_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_8_4_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_8_4_2  (
            .in0(N__36634),
            .in1(_gnd_net_),
            .in2(N__25695),
            .in3(N__26741),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49951),
            .ce(N__31223),
            .sr(N__49349));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_8_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_8_4_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_8_4_4  (
            .in0(N__25691),
            .in1(N__27982),
            .in2(N__25682),
            .in3(N__28000),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_8_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_8_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_8_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_8_4_7  (
            .in0(N__28344),
            .in1(N__28371),
            .in2(_gnd_net_),
            .in3(N__36635),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49951),
            .ce(N__31223),
            .sr(N__49349));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_5_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_5_0  (
            .in0(N__25845),
            .in1(N__27947),
            .in2(N__25614),
            .in3(N__27965),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_5_2  (
            .in0(N__26587),
            .in1(N__25628),
            .in2(_gnd_net_),
            .in3(N__36638),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_8_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_8_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_8_5_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_8_5_3  (
            .in0(N__36640),
            .in1(_gnd_net_),
            .in2(N__25617),
            .in3(N__26588),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49947),
            .ce(N__31211),
            .sr(N__49358));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_8_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_8_5_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_8_5_4  (
            .in0(N__25844),
            .in1(N__27946),
            .in2(N__25613),
            .in3(N__27964),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_8_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_8_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_8_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_8_5_5  (
            .in0(N__36639),
            .in1(N__28632),
            .in2(_gnd_net_),
            .in3(N__28611),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49947),
            .ce(N__31211),
            .sr(N__49358));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_8_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_8_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_8_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_8_5_7  (
            .in0(N__36641),
            .in1(N__31004),
            .in2(_gnd_net_),
            .in3(N__30977),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49947),
            .ce(N__31211),
            .sr(N__49358));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_6_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_6_0  (
            .in0(N__28244),
            .in1(N__28265),
            .in2(N__25803),
            .in3(N__25791),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_8_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_8_6_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_8_6_1  (
            .in0(N__25790),
            .in1(N__28243),
            .in2(N__28269),
            .in3(N__25799),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_8_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_8_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_8_6_2  (
            .in0(N__28916),
            .in1(N__28877),
            .in2(_gnd_net_),
            .in3(N__36542),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_8_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_8_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_8_6_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_8_6_3  (
            .in0(N__36544),
            .in1(_gnd_net_),
            .in2(N__25806),
            .in3(N__28917),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(N__31265),
            .sr(N__49365));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_8_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_8_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_8_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_8_6_5  (
            .in0(N__36543),
            .in1(N__30632),
            .in2(_gnd_net_),
            .in3(N__30606),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(N__31265),
            .sr(N__49365));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_8_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_8_6_7 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_8_6_7  (
            .in0(N__25775),
            .in1(N__28189),
            .in2(N__25764),
            .in3(N__28216),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_8_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_8_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_8_7_0  (
            .in0(N__25986),
            .in1(N__30075),
            .in2(N__28542),
            .in3(N__30145),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_8_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_8_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_8_7_3  (
            .in0(N__30076),
            .in1(N__30103),
            .in2(_gnd_net_),
            .in3(N__36597),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(N__31201),
            .sr(N__49371));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_8_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_8_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_8_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_8_7_7  (
            .in0(N__28563),
            .in1(N__28540),
            .in2(_gnd_net_),
            .in3(N__36598),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(N__31201),
            .sr(N__49371));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_0  (
            .in0(N__26578),
            .in1(N__30744),
            .in2(N__30605),
            .in3(N__30885),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_8_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_8_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_8_8_4  (
            .in0(N__26676),
            .in1(N__26731),
            .in2(N__28610),
            .in3(N__28841),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_8_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_8_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_8_8_6  (
            .in0(N__28865),
            .in1(N__28842),
            .in2(_gnd_net_),
            .in3(N__36472),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49915),
            .ce(N__31254),
            .sr(N__49375));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_9_0  (
            .in0(N__36417),
            .in1(N__25875),
            .in2(_gnd_net_),
            .in3(N__26677),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_8_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_8_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_8_9_1  (
            .in0(N__26379),
            .in1(N__31576),
            .in2(N__30264),
            .in3(N__32470),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_8_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_8_9_2 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_8_9_2  (
            .in0(N__36414),
            .in1(N__28798),
            .in2(N__28775),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_8_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_8_9_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_8_9_3  (
            .in0(N__25857),
            .in1(N__30213),
            .in2(N__25941),
            .in3(N__28423),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_8_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_8_9_4 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_8_9_4  (
            .in0(N__28290),
            .in1(N__25947),
            .in2(N__25848),
            .in3(N__28965),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_8_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_8_9_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__28631),
            .in2(N__25953),
            .in3(N__28605),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_9_6  (
            .in0(N__36415),
            .in1(N__28562),
            .in2(_gnd_net_),
            .in3(N__28541),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_8_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_8_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_8_9_7  (
            .in0(N__28966),
            .in1(N__28937),
            .in2(_gnd_net_),
            .in3(N__36416),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_10_0  (
            .in0(N__30631),
            .in1(N__30597),
            .in2(_gnd_net_),
            .in3(N__36406),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_10_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_10_1  (
            .in0(N__31391),
            .in1(N__32662),
            .in2(N__28477),
            .in3(N__28362),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_10_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__33057),
            .in2(N__25950),
            .in3(N__28910),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_10_3  (
            .in0(N__36407),
            .in1(N__28343),
            .in2(_gnd_net_),
            .in3(N__28363),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_10_4  (
            .in0(N__28864),
            .in1(N__28840),
            .in2(_gnd_net_),
            .in3(N__36408),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_8_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_8_10_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_8_10_6  (
            .in0(N__26125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30960),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__26210),
            .in2(N__25932),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49879),
            .ce(N__27063),
            .sr(N__49389));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__26186),
            .in2(N__26241),
            .in3(N__26214),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49879),
            .ce(N__27063),
            .sr(N__49389));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__26211),
            .in2(N__26165),
            .in3(N__26190),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49879),
            .ce(N__27063),
            .sr(N__49389));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__26187),
            .in2(N__26105),
            .in3(N__26169),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49879),
            .ce(N__27063),
            .sr(N__49389));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__26075),
            .in2(N__26166),
            .in3(N__26109),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49879),
            .ce(N__27063),
            .sr(N__49389));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__26048),
            .in2(N__26106),
            .in3(N__26082),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49879),
            .ce(N__27063),
            .sr(N__49389));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__26018),
            .in2(N__26079),
            .in3(N__26055),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49879),
            .ce(N__27063),
            .sr(N__49389));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__26492),
            .in2(N__26052),
            .in3(N__26025),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49879),
            .ce(N__27063),
            .sr(N__49389));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__26462),
            .in2(N__26022),
            .in3(N__25956),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49869),
            .ce(N__27062),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__26438),
            .in2(N__26499),
            .in3(N__26469),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49869),
            .ce(N__27062),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__26414),
            .in2(N__26466),
            .in3(N__26442),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49869),
            .ce(N__27062),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__26439),
            .in2(N__26351),
            .in3(N__26418),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49869),
            .ce(N__27062),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__26415),
            .in2(N__26324),
            .in3(N__26355),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49869),
            .ce(N__27062),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__26291),
            .in2(N__26352),
            .in3(N__26328),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49869),
            .ce(N__27062),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__26264),
            .in2(N__26325),
            .in3(N__26298),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49869),
            .ce(N__27062),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__26804),
            .in2(N__26295),
            .in3(N__26271),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49869),
            .ce(N__27062),
            .sr(N__49394));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__26780),
            .in2(N__26268),
            .in3(N__26244),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49859),
            .ce(N__27060),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__26759),
            .in2(N__26808),
            .in3(N__26784),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49859),
            .ce(N__27060),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__26781),
            .in2(N__26709),
            .in3(N__26763),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49859),
            .ce(N__27060),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__26760),
            .in2(N__26642),
            .in3(N__26712),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49859),
            .ce(N__27060),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__26708),
            .in2(N__26612),
            .in3(N__26646),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49859),
            .ce(N__27060),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__26552),
            .in2(N__26643),
            .in3(N__26616),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49859),
            .ce(N__27060),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__26522),
            .in2(N__26613),
            .in3(N__26559),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49859),
            .ce(N__27060),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__27173),
            .in2(N__26556),
            .in3(N__26529),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49859),
            .ce(N__27060),
            .sr(N__49397));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__27131),
            .in2(N__26526),
            .in3(N__26502),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49846),
            .ce(N__27059),
            .sr(N__49402));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__27089),
            .in2(N__27177),
            .in3(N__27153),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49846),
            .ce(N__27059),
            .sr(N__49402));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__27150),
            .in2(N__27135),
            .in3(N__27111),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49846),
            .ce(N__27059),
            .sr(N__49402));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__27108),
            .in2(N__27093),
            .in3(N__27069),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49846),
            .ce(N__27059),
            .sr(N__49402));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27066),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(N__27059),
            .sr(N__49402));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_23_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_23_1 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_23_1  (
            .in0(N__26988),
            .in1(N__26934),
            .in2(N__48730),
            .in3(N__26878),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_24_0  (
            .in0(_gnd_net_),
            .in1(N__26850),
            .in2(N__26859),
            .in3(N__27567),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_8_24_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_24_1  (
            .in0(_gnd_net_),
            .in1(N__26832),
            .in2(N__26844),
            .in3(N__27501),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_24_2  (
            .in0(_gnd_net_),
            .in1(N__26814),
            .in2(N__26826),
            .in3(N__27543),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_24_3  (
            .in0(_gnd_net_),
            .in1(N__27318),
            .in2(N__27327),
            .in3(N__27477),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_24_4  (
            .in0(_gnd_net_),
            .in1(N__27297),
            .in2(N__27312),
            .in3(N__27522),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_24_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_24_5  (
            .in0(N__27426),
            .in1(N__27276),
            .in2(N__27291),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_24_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_24_6  (
            .in0(N__27450),
            .in1(N__27261),
            .in2(N__27270),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_24_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_24_7  (
            .in0(N__27588),
            .in1(N__27246),
            .in2(N__27255),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_25_0  (
            .in0(_gnd_net_),
            .in1(N__27228),
            .in2(N__27237),
            .in3(N__27630),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_8_25_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_25_1  (
            .in0(_gnd_net_),
            .in1(N__27210),
            .in2(N__27222),
            .in3(N__27609),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_8_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_8_25_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_8_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_8_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27204),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49806),
            .ce(),
            .sr(N__49446));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_8_26_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_8_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_8_26_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_8_26_0  (
            .in0(N__27625),
            .in1(N__27604),
            .in2(_gnd_net_),
            .in3(N__27586),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_8_26_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_8_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_8_26_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_8_26_5  (
            .in0(_gnd_net_),
            .in1(N__27562),
            .in2(_gnd_net_),
            .in3(N__27538),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_8_26_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_8_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_8_26_6 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_8_26_6  (
            .in0(N__27520),
            .in1(N__27499),
            .in2(N__27480),
            .in3(N__27475),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_8_26_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_8_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_8_26_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_8_26_7  (
            .in0(N__27456),
            .in1(N__27449),
            .in2(N__27429),
            .in3(N__27425),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_2.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_2 (
            .in0(N__27363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_9_1_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_9_1_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_9_1_2 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_9_1_2  (
            .in0(N__32616),
            .in1(N__30000),
            .in2(N__27788),
            .in3(N__31232),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49955),
            .ce(),
            .sr(N__49316));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_2_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_2_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_2_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_9_2_1  (
            .in0(N__30303),
            .in1(_gnd_net_),
            .in2(N__36721),
            .in3(N__30271),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49954),
            .ce(N__31250),
            .sr(N__49324));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_2_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_2_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_2_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_9_2_4  (
            .in0(N__28437),
            .in1(N__36704),
            .in2(_gnd_net_),
            .in3(N__28395),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49954),
            .ce(N__31250),
            .sr(N__49324));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_2_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_2_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_2_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_9_2_5  (
            .in0(N__32639),
            .in1(_gnd_net_),
            .in2(N__36722),
            .in3(N__32691),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49954),
            .ce(N__31250),
            .sr(N__49324));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_9_3_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_9_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(N__29718),
            .in2(N__27789),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_9_3_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_9_3_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_9_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_9_3_1  (
            .in0(N__31117),
            .in1(N__27761),
            .in2(_gnd_net_),
            .in3(N__27747),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49952),
            .ce(),
            .sr(N__49332));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_9_3_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_9_3_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_9_3_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_9_3_2  (
            .in0(N__31121),
            .in1(N__27743),
            .in2(N__29985),
            .in3(N__27729),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49952),
            .ce(),
            .sr(N__49332));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_9_3_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_9_3_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_9_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_9_3_3  (
            .in0(N__31118),
            .in1(N__27725),
            .in2(_gnd_net_),
            .in3(N__27711),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49952),
            .ce(),
            .sr(N__49332));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_9_3_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_9_3_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_9_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_9_3_4  (
            .in0(N__31122),
            .in1(N__27707),
            .in2(_gnd_net_),
            .in3(N__27693),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49952),
            .ce(),
            .sr(N__49332));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_9_3_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_9_3_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_9_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_9_3_5  (
            .in0(N__31119),
            .in1(N__27689),
            .in2(_gnd_net_),
            .in3(N__27675),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49952),
            .ce(),
            .sr(N__49332));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_3_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_3_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_3_6  (
            .in0(N__31123),
            .in1(N__27668),
            .in2(_gnd_net_),
            .in3(N__27654),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49952),
            .ce(),
            .sr(N__49332));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_3_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_3_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_3_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_3_7  (
            .in0(N__31120),
            .in1(N__27650),
            .in2(_gnd_net_),
            .in3(N__27633),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49952),
            .ce(),
            .sr(N__49332));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_4_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_4_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_4_0  (
            .in0(N__31219),
            .in1(N__27929),
            .in2(_gnd_net_),
            .in3(N__27915),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49948),
            .ce(),
            .sr(N__49341));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_9_4_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_9_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_9_4_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_9_4_1  (
            .in0(N__31212),
            .in1(N__27911),
            .in2(_gnd_net_),
            .in3(N__27897),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49948),
            .ce(),
            .sr(N__49341));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_9_4_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_9_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_9_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_9_4_2  (
            .in0(N__31216),
            .in1(N__27893),
            .in2(_gnd_net_),
            .in3(N__27879),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49948),
            .ce(),
            .sr(N__49341));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_4_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_4_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_4_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_4_3  (
            .in0(N__31213),
            .in1(N__27875),
            .in2(_gnd_net_),
            .in3(N__27861),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49948),
            .ce(),
            .sr(N__49341));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_9_4_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_9_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_9_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_9_4_4  (
            .in0(N__31217),
            .in1(N__27854),
            .in2(_gnd_net_),
            .in3(N__27840),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49948),
            .ce(),
            .sr(N__49341));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_9_4_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_9_4_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_9_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_9_4_5  (
            .in0(N__31214),
            .in1(N__27833),
            .in2(_gnd_net_),
            .in3(N__27819),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49948),
            .ce(),
            .sr(N__49341));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_9_4_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_9_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_9_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_9_4_6  (
            .in0(N__31218),
            .in1(N__27815),
            .in2(_gnd_net_),
            .in3(N__27801),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49948),
            .ce(),
            .sr(N__49341));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_9_4_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_9_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_9_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_9_4_7  (
            .in0(N__31215),
            .in1(N__29939),
            .in2(_gnd_net_),
            .in3(N__27798),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49948),
            .ce(),
            .sr(N__49341));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_9_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_9_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_9_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_9_5_0  (
            .in0(N__31224),
            .in1(N__29921),
            .in2(_gnd_net_),
            .in3(N__28113),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49350));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_9_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_9_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_9_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_9_5_1  (
            .in0(N__31228),
            .in1(N__28102),
            .in2(_gnd_net_),
            .in3(N__28080),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49350));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_9_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_9_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_9_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_9_5_2  (
            .in0(N__31225),
            .in1(N__28075),
            .in2(_gnd_net_),
            .in3(N__28053),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49350));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_9_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_9_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_9_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_9_5_3  (
            .in0(N__31229),
            .in1(N__28048),
            .in2(_gnd_net_),
            .in3(N__28032),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49350));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_9_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_9_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_9_5_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_9_5_4  (
            .in0(N__31226),
            .in1(_gnd_net_),
            .in2(N__28028),
            .in3(N__28005),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49350));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_9_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_9_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_9_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_9_5_5  (
            .in0(N__31230),
            .in1(N__28002),
            .in2(_gnd_net_),
            .in3(N__27987),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49350));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_9_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_9_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_9_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_9_5_6  (
            .in0(N__31227),
            .in1(N__27984),
            .in2(_gnd_net_),
            .in3(N__27969),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49350));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_9_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_9_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_9_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_9_5_7  (
            .in0(N__31231),
            .in1(N__27966),
            .in2(_gnd_net_),
            .in3(N__27951),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49938),
            .ce(),
            .sr(N__49350));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_9_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_9_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_9_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_9_6_0  (
            .in0(N__31233),
            .in1(N__27948),
            .in2(_gnd_net_),
            .in3(N__27933),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49928),
            .ce(),
            .sr(N__49359));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_9_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_9_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_9_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_9_6_1  (
            .in0(N__31237),
            .in1(N__28264),
            .in2(_gnd_net_),
            .in3(N__28248),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49928),
            .ce(),
            .sr(N__49359));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_9_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_9_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_9_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_9_6_2  (
            .in0(N__31234),
            .in1(N__28245),
            .in2(_gnd_net_),
            .in3(N__28230),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49928),
            .ce(),
            .sr(N__49359));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_9_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_9_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_9_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_9_6_3  (
            .in0(N__31238),
            .in1(N__28145),
            .in2(_gnd_net_),
            .in3(N__28227),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49928),
            .ce(),
            .sr(N__49359));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_9_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_9_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_9_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_9_6_4  (
            .in0(N__31235),
            .in1(N__28161),
            .in2(_gnd_net_),
            .in3(N__28224),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49928),
            .ce(),
            .sr(N__49359));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_9_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_9_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_9_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_9_6_5  (
            .in0(N__31239),
            .in1(N__28220),
            .in2(_gnd_net_),
            .in3(N__28200),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49928),
            .ce(),
            .sr(N__49359));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_9_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_9_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_9_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_9_6_6  (
            .in0(N__31236),
            .in1(N__28193),
            .in2(_gnd_net_),
            .in3(N__28197),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49359));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_7_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_7_0  (
            .in0(N__28160),
            .in1(N__28141),
            .in2(N__28323),
            .in3(N__29874),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_7_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_7_1  (
            .in0(N__29873),
            .in1(N__28159),
            .in2(N__28146),
            .in3(N__28319),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_9_7_3  (
            .in0(N__30769),
            .in1(N__30753),
            .in2(_gnd_net_),
            .in3(N__36682),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(N__31264),
            .sr(N__49366));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_8_0  (
            .in0(N__36413),
            .in1(N__30105),
            .in2(_gnd_net_),
            .in3(N__30083),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_9_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_9_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_9_8_1  (
            .in0(N__30773),
            .in1(N__30752),
            .in2(_gnd_net_),
            .in3(N__36409),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2  (
            .in0(N__28768),
            .in1(N__31348),
            .in2(N__33204),
            .in3(N__36762),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_3  (
            .in0(N__28311),
            .in1(N__28305),
            .in2(N__28299),
            .in3(N__28296),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_8_4  (
            .in0(N__36412),
            .in1(N__28430),
            .in2(_gnd_net_),
            .in3(N__28393),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_9_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_9_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_9_8_5  (
            .in0(N__31000),
            .in1(N__30970),
            .in2(_gnd_net_),
            .in3(N__36410),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_8_7  (
            .in0(N__33067),
            .in1(N__33026),
            .in2(_gnd_net_),
            .in3(N__36411),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_9_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_9_0  (
            .in0(N__31751),
            .in1(N__28280),
            .in2(N__31728),
            .in3(N__28572),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_9_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_9_1  (
            .in0(N__28571),
            .in1(N__31727),
            .in2(N__28284),
            .in3(N__31752),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_9_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_9_9_2  (
            .in0(N__36467),
            .in1(N__28627),
            .in2(_gnd_net_),
            .in3(N__28609),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49893),
            .ce(N__33335),
            .sr(N__49376));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_9_9_7  (
            .in0(N__28558),
            .in1(N__28536),
            .in2(_gnd_net_),
            .in3(N__36468),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49893),
            .ce(N__33335),
            .sr(N__49376));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_10_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_10_0  (
            .in0(N__31841),
            .in1(N__28811),
            .in2(N__31821),
            .in3(N__28446),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_9_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_9_10_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_9_10_1  (
            .in0(N__28445),
            .in1(N__31820),
            .in2(N__28815),
            .in3(N__31842),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_9_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_9_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_9_10_4  (
            .in0(N__28509),
            .in1(N__28482),
            .in2(_gnd_net_),
            .in3(N__36473),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49880),
            .ce(N__33337),
            .sr(N__49381));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_9_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_9_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_9_11_3  (
            .in0(N__33155),
            .in1(N__33201),
            .in2(_gnd_net_),
            .in3(N__36560),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(N__33340),
            .sr(N__49386));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_9_11_4  (
            .in0(N__36672),
            .in1(N__28422),
            .in2(_gnd_net_),
            .in3(N__28394),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(N__33340),
            .sr(N__49386));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_9_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_9_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_9_11_5  (
            .in0(N__28364),
            .in1(N__28339),
            .in2(_gnd_net_),
            .in3(N__36561),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(N__33340),
            .sr(N__49386));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_9_11_7  (
            .in0(N__31314),
            .in1(N__31338),
            .in2(_gnd_net_),
            .in3(N__36559),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49870),
            .ce(N__33340),
            .sr(N__49386));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_9_12_1  (
            .in0(N__28973),
            .in1(N__28938),
            .in2(_gnd_net_),
            .in3(N__36558),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(N__33341),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_9_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_9_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_9_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_9_12_4  (
            .in0(N__36555),
            .in1(N__28909),
            .in2(_gnd_net_),
            .in3(N__28884),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(N__33341),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_9_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_9_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_9_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_9_12_5  (
            .in0(N__28866),
            .in1(N__28834),
            .in2(_gnd_net_),
            .in3(N__36557),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(N__33341),
            .sr(N__49390));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_9_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_9_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_9_12_7  (
            .in0(N__28800),
            .in1(N__28758),
            .in2(_gnd_net_),
            .in3(N__36556),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(N__33341),
            .sr(N__49390));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_13_0  (
            .in0(N__31899),
            .in1(N__28740),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_9_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_9_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_9_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__32127),
            .in2(_gnd_net_),
            .in3(N__28698),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__49847),
            .ce(),
            .sr(N__49395));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_9_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_9_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_9_13_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32115),
            .in3(N__28668),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__49847),
            .ce(),
            .sr(N__49395));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_9_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_9_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_9_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__32100),
            .in2(_gnd_net_),
            .in3(N__28635),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__49847),
            .ce(),
            .sr(N__49395));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_9_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_9_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_9_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__32088),
            .in2(_gnd_net_),
            .in3(N__29217),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__49847),
            .ce(),
            .sr(N__49395));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_9_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_9_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_9_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32076),
            .in3(N__29196),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__49847),
            .ce(),
            .sr(N__49395));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_9_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_9_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_9_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__32061),
            .in2(_gnd_net_),
            .in3(N__29172),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__49847),
            .ce(),
            .sr(N__49395));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_9_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_9_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_9_13_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32049),
            .in3(N__29142),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__49847),
            .ce(),
            .sr(N__49395));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_9_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_9_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_9_14_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32034),
            .in3(N__29109),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__49837),
            .ce(),
            .sr(N__49398));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_9_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_9_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__32019),
            .in2(_gnd_net_),
            .in3(N__29079),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__49837),
            .ce(),
            .sr(N__49398));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_9_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_9_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_9_14_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32235),
            .in3(N__29046),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__49837),
            .ce(),
            .sr(N__49398));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_9_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_9_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_9_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__32220),
            .in2(_gnd_net_),
            .in3(N__29013),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__49837),
            .ce(),
            .sr(N__49398));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_9_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_9_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__32208),
            .in2(_gnd_net_),
            .in3(N__28977),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__49837),
            .ce(),
            .sr(N__49398));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_9_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_9_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_9_14_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32196),
            .in3(N__29448),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__49837),
            .ce(),
            .sr(N__49398));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_9_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_9_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_9_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__32181),
            .in2(_gnd_net_),
            .in3(N__29418),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__49837),
            .ce(),
            .sr(N__49398));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_9_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_9_14_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32169),
            .in3(N__29394),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__49837),
            .ce(),
            .sr(N__49398));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_9_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_9_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_9_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__32154),
            .in2(_gnd_net_),
            .in3(N__29361),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__49828),
            .ce(),
            .sr(N__49403));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_9_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_9_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_9_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32142),
            .in3(N__29337),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__49828),
            .ce(),
            .sr(N__49403));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_9_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_9_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__32340),
            .in2(_gnd_net_),
            .in3(N__29307),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__49828),
            .ce(),
            .sr(N__49403));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_9_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_9_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_9_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__32328),
            .in2(_gnd_net_),
            .in3(N__29274),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__49828),
            .ce(),
            .sr(N__49403));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_9_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_9_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_9_15_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32316),
            .in3(N__29247),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__49828),
            .ce(),
            .sr(N__49403));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_9_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_9_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_9_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__32301),
            .in2(_gnd_net_),
            .in3(N__29688),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__49828),
            .ce(),
            .sr(N__49403));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_9_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_9_15_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32289),
            .in3(N__29658),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__49828),
            .ce(),
            .sr(N__49403));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_9_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_9_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_9_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32274),
            .in3(N__29631),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__49828),
            .ce(),
            .sr(N__49403));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_9_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_9_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_9_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__32259),
            .in2(_gnd_net_),
            .in3(N__29601),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__49822),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_9_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_9_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_9_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__32247),
            .in2(_gnd_net_),
            .in3(N__29568),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__49822),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_9_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_9_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_9_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__32448),
            .in2(_gnd_net_),
            .in3(N__29535),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .clk(N__49822),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_9_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_9_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_9_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_27_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__32436),
            .in2(_gnd_net_),
            .in3(N__29502),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .clk(N__49822),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_9_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_9_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_9_16_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_28_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32424),
            .in3(N__29472),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .clk(N__49822),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_9_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_9_16_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_29_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32409),
            .in3(N__29841),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .clk(N__49822),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_9_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_9_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_9_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_30_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__30717),
            .in2(_gnd_net_),
            .in3(N__29811),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ),
            .clk(N__49822),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_9_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_9_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_9_16_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_31_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__32391),
            .in2(_gnd_net_),
            .in3(N__29808),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49822),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29805),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49814),
            .ce(),
            .sr(N__49426));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29787),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49808),
            .ce(),
            .sr(N__49437));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_1_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_1_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_10_1_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_10_1_6  (
            .in0(N__31376),
            .in1(N__31419),
            .in2(_gnd_net_),
            .in3(N__36702),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49953),
            .ce(N__31256),
            .sr(N__49302));
    defparam \phase_controller_inst1.stoper_tr.running_LC_10_3_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_10_3_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_10_3_3 .LUT_INIT=16'b1100010011101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_10_3_3  (
            .in0(N__32605),
            .in1(N__31431),
            .in2(N__32583),
            .in3(N__32535),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49939),
            .ce(),
            .sr(N__49317));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_10_3_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_10_3_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_10_3_5  (
            .in0(_gnd_net_),
            .in1(N__32534),
            .in2(_gnd_net_),
            .in3(N__32575),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_10_3_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_10_3_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_10_3_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_10_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29721),
            .in3(N__32603),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_10_3_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_10_3_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_10_3_7  (
            .in0(N__32604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29996),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_10_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_10_4_2  (
            .in0(N__30121),
            .in1(N__30162),
            .in2(_gnd_net_),
            .in3(N__36712),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49929),
            .ce(N__31199),
            .sr(N__49325));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_10_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_10_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_10_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_10_4_4  (
            .in0(N__32506),
            .in1(N__32486),
            .in2(_gnd_net_),
            .in3(N__36711),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49929),
            .ce(N__31199),
            .sr(N__49325));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_5_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_5_0  (
            .in0(N__29917),
            .in1(N__29886),
            .in2(N__29940),
            .in3(N__29949),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_5_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_5_1  (
            .in0(N__29948),
            .in1(N__29938),
            .in2(N__29922),
            .in3(N__29885),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_5_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_5_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_5_6  (
            .in0(N__36631),
            .in1(N__30125),
            .in2(_gnd_net_),
            .in3(N__30154),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_5_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_5_7  (
            .in0(N__30298),
            .in1(N__36630),
            .in2(_gnd_net_),
            .in3(N__30278),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_10_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_10_6_3  (
            .in0(N__36237),
            .in1(N__36773),
            .in2(_gnd_net_),
            .in3(N__36679),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49906),
            .ce(N__31266),
            .sr(N__49342));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_10_6_7  (
            .in0(N__33072),
            .in1(N__33022),
            .in2(_gnd_net_),
            .in3(N__36680),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49906),
            .ce(N__31266),
            .sr(N__49342));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_10_7_0  (
            .in0(N__36673),
            .in1(N__30299),
            .in2(_gnd_net_),
            .in3(N__30279),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49895),
            .ce(N__33333),
            .sr(N__49351));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_10_7_1  (
            .in0(N__30227),
            .in1(N__30189),
            .in2(_gnd_net_),
            .in3(N__36677),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49895),
            .ce(N__33333),
            .sr(N__49351));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_10_7_2  (
            .in0(N__36674),
            .in1(N__32646),
            .in2(_gnd_net_),
            .in3(N__32683),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49895),
            .ce(N__33333),
            .sr(N__49351));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_10_7_3  (
            .in0(N__30161),
            .in1(N__30126),
            .in2(_gnd_net_),
            .in3(N__36678),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49895),
            .ce(N__33333),
            .sr(N__49351));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_10_7_4  (
            .in0(N__36675),
            .in1(N__31380),
            .in2(_gnd_net_),
            .in3(N__31418),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49895),
            .ce(N__33333),
            .sr(N__49351));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_10_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_10_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_10_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_10_7_5  (
            .in0(N__30104),
            .in1(N__30087),
            .in2(_gnd_net_),
            .in3(N__36676),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49895),
            .ce(N__33333),
            .sr(N__49351));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_10_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_10_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__30039),
            .in2(N__30048),
            .in3(N__32770),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_10_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_10_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__30021),
            .in2(N__30033),
            .in3(N__31535),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_10_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_10_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__30006),
            .in2(N__30015),
            .in3(N__31520),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_10_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_10_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__30441),
            .in2(N__30432),
            .in3(N__31505),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_10_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_10_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__30423),
            .in2(N__30417),
            .in3(N__31490),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_10_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_10_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__30405),
            .in2(N__30396),
            .in3(N__31475),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_10_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_10_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__30387),
            .in2(N__30375),
            .in3(N__31460),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_10_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_10_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_10_8_7  (
            .in0(N__31445),
            .in1(N__30945),
            .in2(N__30366),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_10_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_10_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__30357),
            .in2(N__30348),
            .in3(N__31700),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_10_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_10_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__30339),
            .in2(N__30330),
            .in3(N__31685),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_10_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_10_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__30321),
            .in2(N__30312),
            .in3(N__31670),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_10_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_10_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__30534),
            .in2(N__30543),
            .in3(N__31655),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_10_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_10_9_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_10_9_4  (
            .in0(N__31640),
            .in1(N__30528),
            .in2(N__30519),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_10_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_10_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__30510),
            .in2(N__31548),
            .in3(N__31625),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_10_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_10_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__30504),
            .in2(N__30489),
            .in3(N__31610),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_10_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_10_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__33099),
            .in2(N__32940),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_10_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_10_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__30816),
            .in2(N__30849),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_10_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_10_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__30480),
            .in2(N__30474),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_10_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_10_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__30462),
            .in2(N__30453),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_10_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_10_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__30678),
            .in2(N__30672),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_10_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_10_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__30639),
            .in2(N__30660),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_10_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_10_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__33222),
            .in2(N__33087),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_10_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_10_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__30927),
            .in2(N__30552),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30663),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_11_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_11_0  (
            .in0(N__32005),
            .in1(N__31988),
            .in2(N__30651),
            .in3(N__30561),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_10_11_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_10_11_1  (
            .in0(N__30560),
            .in1(N__32006),
            .in2(N__31989),
            .in3(N__30650),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_10_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_10_11_2  (
            .in0(N__30633),
            .in1(N__30604),
            .in2(_gnd_net_),
            .in3(N__36671),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49849),
            .ce(N__33336),
            .sr(N__49377));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_10_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_10_11_5 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_10_11_5  (
            .in0(N__30857),
            .in1(N__31934),
            .in2(N__30939),
            .in3(N__31957),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_6 .LUT_INIT=16'b0010101100100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_6  (
            .in0(N__31933),
            .in1(N__30938),
            .in2(N__31959),
            .in3(N__30858),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_10_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_10_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_10_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_10_11_7  (
            .in0(N__36670),
            .in1(N__30921),
            .in2(_gnd_net_),
            .in3(N__30894),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49849),
            .ce(N__33336),
            .sr(N__49377));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_12_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_12_0  (
            .in0(N__31862),
            .in1(N__30824),
            .in2(N__31887),
            .in3(N__30837),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_12_1 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_12_1  (
            .in0(N__30836),
            .in1(N__31886),
            .in2(N__30828),
            .in3(N__31863),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_10_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__31919),
            .in2(_gnd_net_),
            .in3(N__37830),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(N__49387));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_10_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_10_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_10_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_10_14_5  (
            .in0(N__30777),
            .in1(N__30751),
            .in2(_gnd_net_),
            .in3(N__36714),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49823),
            .ce(N__33342),
            .sr(N__49391));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32387),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_0 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_0  (
            .in0(N__48891),
            .in1(N__30711),
            .in2(N__48729),
            .in3(N__48932),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_3_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_3_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_3_1  (
            .in0(N__32526),
            .in1(N__31430),
            .in2(_gnd_net_),
            .in3(N__32550),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_11_3_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_11_3_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_11_3_6  (
            .in0(N__32551),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32527),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_11_4_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_11_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_11_4_2  (
            .in0(N__31375),
            .in1(N__31414),
            .in2(_gnd_net_),
            .in3(N__36687),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_5_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_5_3  (
            .in0(N__32508),
            .in1(N__32485),
            .in2(_gnd_net_),
            .in3(N__36688),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_5_7 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_5_7  (
            .in0(N__32887),
            .in1(N__33724),
            .in2(N__38322),
            .in3(N__32847),
            .lcout(\phase_controller_inst2.N_54_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_11_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_11_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_11_6_1  (
            .in0(N__31306),
            .in1(N__31355),
            .in2(_gnd_net_),
            .in3(N__36689),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_11_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_11_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_11_6_5  (
            .in0(N__31591),
            .in1(N__31559),
            .in2(_gnd_net_),
            .in3(N__36690),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_11_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_11_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_11_6_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_11_6_6  (
            .in0(N__36691),
            .in1(_gnd_net_),
            .in2(N__31284),
            .in3(N__31592),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49896),
            .ce(N__31263),
            .sr(N__49333));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_11_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_11_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_11_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_11_7_0  (
            .in0(N__31005),
            .in1(N__30978),
            .in2(_gnd_net_),
            .in3(N__36701),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49881),
            .ce(N__33332),
            .sr(N__49343));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_11_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_11_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_11_7_6  (
            .in0(N__31593),
            .in1(N__31560),
            .in2(_gnd_net_),
            .in3(N__36700),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49881),
            .ce(N__33332),
            .sr(N__49343));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__32709),
            .in2(N__32771),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_11_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_11_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_11_8_1  (
            .in0(N__33668),
            .in1(N__31536),
            .in2(_gnd_net_),
            .in3(N__31524),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49872),
            .ce(),
            .sr(N__49352));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_11_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_11_8_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_11_8_2  (
            .in0(N__33676),
            .in1(N__31521),
            .in2(N__33132),
            .in3(N__31509),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49872),
            .ce(),
            .sr(N__49352));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_11_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_11_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_11_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_11_8_3  (
            .in0(N__33669),
            .in1(N__31506),
            .in2(_gnd_net_),
            .in3(N__31494),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49872),
            .ce(),
            .sr(N__49352));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_11_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_11_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_11_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_11_8_4  (
            .in0(N__33677),
            .in1(N__31491),
            .in2(_gnd_net_),
            .in3(N__31479),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49872),
            .ce(),
            .sr(N__49352));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_11_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_11_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_11_8_5  (
            .in0(N__33670),
            .in1(N__31476),
            .in2(_gnd_net_),
            .in3(N__31464),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49872),
            .ce(),
            .sr(N__49352));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_11_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_11_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_11_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_11_8_6  (
            .in0(N__33678),
            .in1(N__31461),
            .in2(_gnd_net_),
            .in3(N__31449),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49872),
            .ce(),
            .sr(N__49352));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_11_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_11_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_11_8_7  (
            .in0(N__33671),
            .in1(N__31446),
            .in2(_gnd_net_),
            .in3(N__31434),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49872),
            .ce(),
            .sr(N__49352));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_11_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_11_9_0  (
            .in0(N__33675),
            .in1(N__31701),
            .in2(_gnd_net_),
            .in3(N__31689),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49862),
            .ce(),
            .sr(N__49360));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_11_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_11_9_1  (
            .in0(N__33679),
            .in1(N__31686),
            .in2(_gnd_net_),
            .in3(N__31674),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49862),
            .ce(),
            .sr(N__49360));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_11_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_11_9_2  (
            .in0(N__33672),
            .in1(N__31671),
            .in2(_gnd_net_),
            .in3(N__31659),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49862),
            .ce(),
            .sr(N__49360));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_11_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_11_9_3  (
            .in0(N__33680),
            .in1(N__31656),
            .in2(_gnd_net_),
            .in3(N__31644),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49862),
            .ce(),
            .sr(N__49360));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_11_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_11_9_4  (
            .in0(N__33673),
            .in1(N__31641),
            .in2(_gnd_net_),
            .in3(N__31629),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49862),
            .ce(),
            .sr(N__49360));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_11_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_11_9_5  (
            .in0(N__33681),
            .in1(N__31626),
            .in2(_gnd_net_),
            .in3(N__31614),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49862),
            .ce(),
            .sr(N__49360));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_11_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_11_9_6  (
            .in0(N__33674),
            .in1(N__31611),
            .in2(_gnd_net_),
            .in3(N__31599),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49862),
            .ce(),
            .sr(N__49360));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_11_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_11_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_11_9_7  (
            .in0(N__33682),
            .in1(N__32962),
            .in2(_gnd_net_),
            .in3(N__31596),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49862),
            .ce(),
            .sr(N__49360));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_11_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_11_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_11_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_11_10_0  (
            .in0(N__33692),
            .in1(N__33000),
            .in2(_gnd_net_),
            .in3(N__31890),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49850),
            .ce(),
            .sr(N__49367));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_11_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_11_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_11_10_1  (
            .in0(N__33696),
            .in1(N__31882),
            .in2(_gnd_net_),
            .in3(N__31866),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49850),
            .ce(),
            .sr(N__49367));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_11_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_11_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_11_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_11_10_2  (
            .in0(N__33693),
            .in1(N__31861),
            .in2(_gnd_net_),
            .in3(N__31845),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49850),
            .ce(),
            .sr(N__49367));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_11_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_11_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_11_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_11_10_3  (
            .in0(N__33697),
            .in1(N__31840),
            .in2(_gnd_net_),
            .in3(N__31824),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49850),
            .ce(),
            .sr(N__49367));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_11_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_11_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_11_10_4  (
            .in0(N__33694),
            .in1(N__31816),
            .in2(_gnd_net_),
            .in3(N__31800),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49850),
            .ce(),
            .sr(N__49367));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_11_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_11_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_11_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_11_10_5  (
            .in0(N__33698),
            .in1(N__31792),
            .in2(_gnd_net_),
            .in3(N__31776),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49850),
            .ce(),
            .sr(N__49367));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_11_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_11_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_11_10_6  (
            .in0(N__33695),
            .in1(N__31771),
            .in2(_gnd_net_),
            .in3(N__31755),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49850),
            .ce(),
            .sr(N__49367));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_11_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_11_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_11_10_7  (
            .in0(N__33699),
            .in1(N__31745),
            .in2(_gnd_net_),
            .in3(N__31731),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49850),
            .ce(),
            .sr(N__49367));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_11_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_11_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_11_11_0  (
            .in0(N__33689),
            .in1(N__31718),
            .in2(_gnd_net_),
            .in3(N__31704),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49839),
            .ce(),
            .sr(N__49372));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_11_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_11_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_11_11_1  (
            .in0(N__33685),
            .in1(N__32007),
            .in2(_gnd_net_),
            .in3(N__31992),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49839),
            .ce(),
            .sr(N__49372));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_11_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_11_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_11_11_2  (
            .in0(N__33690),
            .in1(N__31984),
            .in2(_gnd_net_),
            .in3(N__31968),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49839),
            .ce(),
            .sr(N__49372));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_11_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_11_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_11_11_3  (
            .in0(N__33686),
            .in1(N__33240),
            .in2(_gnd_net_),
            .in3(N__31965),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49839),
            .ce(),
            .sr(N__49372));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_11_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_11_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_11_11_4  (
            .in0(N__33691),
            .in1(N__33282),
            .in2(_gnd_net_),
            .in3(N__31962),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49839),
            .ce(),
            .sr(N__49372));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_11_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_11_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_11_11_5  (
            .in0(N__33687),
            .in1(N__31958),
            .in2(_gnd_net_),
            .in3(N__31941),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49839),
            .ce(),
            .sr(N__49372));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_11_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_11_11_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_11_11_6  (
            .in0(N__31935),
            .in1(N__33688),
            .in2(_gnd_net_),
            .in3(N__31938),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49839),
            .ce(),
            .sr(N__49372));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38489),
            .lcout(\current_shift_inst.N_1263_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__37829),
            .in2(N__31920),
            .in3(N__31918),
            .lcout(\current_shift_inst.control_input_1 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_13_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__37353),
            .in2(_gnd_net_),
            .in3(N__32118),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_13_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__33300),
            .in2(_gnd_net_),
            .in3(N__32103),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_13_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__38022),
            .in2(_gnd_net_),
            .in3(N__32091),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_13_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__38145),
            .in2(_gnd_net_),
            .in3(N__32079),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_13_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__37860),
            .in2(_gnd_net_),
            .in3(N__32064),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__33210),
            .in2(_gnd_net_),
            .in3(N__32052),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_13_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__38100),
            .in2(_gnd_net_),
            .in3(N__32037),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_14_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__38052),
            .in2(_gnd_net_),
            .in3(N__32022),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_14_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__33384),
            .in2(_gnd_net_),
            .in3(N__32010),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__33411),
            .in2(_gnd_net_),
            .in3(N__32223),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_14_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__33366),
            .in2(_gnd_net_),
            .in3(N__32211),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_14_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__33378),
            .in2(_gnd_net_),
            .in3(N__32199),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_14_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__33372),
            .in2(_gnd_net_),
            .in3(N__32184),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_12 ),
            .carryout(\current_shift_inst.control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_14_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__33441),
            .in2(_gnd_net_),
            .in3(N__32172),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_13 ),
            .carryout(\current_shift_inst.control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__33360),
            .in2(_gnd_net_),
            .in3(N__32157),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_14 ),
            .carryout(\current_shift_inst.control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_15_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__33435),
            .in2(_gnd_net_),
            .in3(N__32145),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\current_shift_inst.control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_15_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__32364),
            .in2(_gnd_net_),
            .in3(N__32130),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_16 ),
            .carryout(\current_shift_inst.control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__33429),
            .in2(_gnd_net_),
            .in3(N__32331),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_17 ),
            .carryout(\current_shift_inst.control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_15_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__33423),
            .in2(_gnd_net_),
            .in3(N__32319),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_18 ),
            .carryout(\current_shift_inst.control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_15_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__33417),
            .in2(_gnd_net_),
            .in3(N__32304),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_19 ),
            .carryout(\current_shift_inst.control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__36807),
            .in2(_gnd_net_),
            .in3(N__32292),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_20 ),
            .carryout(\current_shift_inst.control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__36105),
            .in2(_gnd_net_),
            .in3(N__32277),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_21 ),
            .carryout(\current_shift_inst.control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_15_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__33402),
            .in2(_gnd_net_),
            .in3(N__32262),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_22 ),
            .carryout(\current_shift_inst.control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_16_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__33396),
            .in2(_gnd_net_),
            .in3(N__32250),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_16_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__33390),
            .in2(_gnd_net_),
            .in3(N__32238),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_24 ),
            .carryout(\current_shift_inst.control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_16_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__32376),
            .in2(_gnd_net_),
            .in3(N__32439),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_25 ),
            .carryout(\current_shift_inst.control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_16_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__33549),
            .in2(_gnd_net_),
            .in3(N__32427),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_26 ),
            .carryout(\current_shift_inst.control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__36048),
            .in2(_gnd_net_),
            .in3(N__32412),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_27 ),
            .carryout(\current_shift_inst.control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_16_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__32370),
            .in2(_gnd_net_),
            .in3(N__32397),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_28 ),
            .carryout(\current_shift_inst.control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__38496),
            .in2(_gnd_net_),
            .in3(N__32394),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_11_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_11_17_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_11_17_5  (
            .in0(N__34659),
            .in1(N__36093),
            .in2(_gnd_net_),
            .in3(N__38497),
            .lcout(\current_shift_inst.control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_11_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_11_17_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_11_17_6  (
            .in0(N__38498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_18_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_18_1  (
            .in0(N__34566),
            .in1(N__35799),
            .in2(_gnd_net_),
            .in3(N__38479),
            .lcout(\current_shift_inst.control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_11_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_11_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_11_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_11_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32865),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49799),
            .ce(),
            .sr(N__49434));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_2_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_2_1  (
            .in0(N__32638),
            .in1(N__32684),
            .in2(_gnd_net_),
            .in3(N__36686),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_12_2_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_12_2_5 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_12_2_5  (
            .in0(N__33469),
            .in1(N__33802),
            .in2(N__33498),
            .in3(N__34887),
            .lcout(\phase_controller_inst1.state_ns_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_3_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_3_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_3_2 .LUT_INIT=16'b1000110010101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_12_3_2  (
            .in0(N__32533),
            .in1(N__33496),
            .in2(N__32615),
            .in3(N__32582),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49917),
            .ce(),
            .sr(N__49303));
    defparam \phase_controller_inst1.start_timer_tr_LC_12_3_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_12_3_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_12_3_5 .LUT_INIT=16'b0111001111110011;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_12_3_5  (
            .in0(N__33495),
            .in1(N__33840),
            .in2(N__32556),
            .in3(N__33473),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49917),
            .ce(),
            .sr(N__49303));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_12_3_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_12_3_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_12_3_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_12_3_7  (
            .in0(N__32555),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49917),
            .ce(),
            .sr(N__49303));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_12_4_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_12_4_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_12_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_12_4_3  (
            .in0(N__32507),
            .in1(N__32490),
            .in2(_gnd_net_),
            .in3(N__36713),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49905),
            .ce(N__33331),
            .sr(N__49310));
    defparam \phase_controller_inst2.start_timer_hc_LC_12_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_12_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_12_5_2 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_12_5_2  (
            .in0(N__33748),
            .in1(N__33707),
            .in2(N__38979),
            .in3(N__32914),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49894),
            .ce(),
            .sr(N__49318));
    defparam \phase_controller_inst2.state_2_LC_12_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_12_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_12_5_3 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_inst2.state_2_LC_12_5_3  (
            .in0(N__32915),
            .in1(N__38321),
            .in2(N__33729),
            .in3(N__33749),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49894),
            .ce(),
            .sr(N__49318));
    defparam \phase_controller_inst2.state_1_LC_12_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_12_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_12_5_4 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst2.state_1_LC_12_5_4  (
            .in0(N__32854),
            .in1(N__33708),
            .in2(_gnd_net_),
            .in3(N__32888),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49894),
            .ce(),
            .sr(N__49318));
    defparam \phase_controller_inst2.state_RNO_0_3_LC_12_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNO_0_3_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNO_0_3_LC_12_6_6 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \phase_controller_inst2.state_RNO_0_3_LC_12_6_6  (
            .in0(N__32922),
            .in1(N__33747),
            .in2(N__32802),
            .in3(N__32827),
            .lcout(\phase_controller_inst2.state_ns_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_12_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_12_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_12_7_2 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst2.state_0_LC_12_7_2  (
            .in0(N__32895),
            .in1(N__32828),
            .in2(N__32801),
            .in3(N__32858),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49871),
            .ce(),
            .sr(N__49334));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_12_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_12_8_0 .LUT_INIT=16'b1000101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_12_8_0  (
            .in0(N__35710),
            .in1(N__32796),
            .in2(N__32745),
            .in3(N__35622),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(N__49344));
    defparam \phase_controller_inst2.start_timer_tr_LC_12_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_12_8_2 .LUT_INIT=16'b0111001111110011;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_12_8_2  (
            .in0(N__32829),
            .in1(N__32811),
            .in2(N__35656),
            .in3(N__32797),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(N__49344));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_8_4 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_8_4  (
            .in0(N__32703),
            .in1(N__35621),
            .in2(N__32772),
            .in3(N__33683),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(),
            .sr(N__49344));
    defparam \phase_controller_inst2.stoper_tr.running_LC_12_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_12_9_3 .LUT_INIT=16'b1101010111001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_12_9_3  (
            .in0(N__35706),
            .in1(N__35678),
            .in2(N__32744),
            .in3(N__35620),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(N__49353));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_12_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_12_9_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__35705),
            .in2(_gnd_net_),
            .in3(N__32737),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32712),
            .in3(N__35618),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35660),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(N__49353));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_12_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_12_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__35619),
            .in2(_gnd_net_),
            .in3(N__32702),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_10_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_10_0  (
            .in0(N__40847),
            .in1(N__40823),
            .in2(N__33111),
            .in3(N__33120),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_10_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_10_1  (
            .in0(N__33119),
            .in1(N__40848),
            .in2(N__40827),
            .in3(N__33107),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_12_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_12_10_2  (
            .in0(N__39696),
            .in1(N__34269),
            .in2(_gnd_net_),
            .in3(N__47075),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49838),
            .ce(N__47153),
            .sr(N__49361));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_12_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_12_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_12_10_3  (
            .in0(N__47074),
            .in1(N__39654),
            .in2(_gnd_net_),
            .in3(N__34250),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49838),
            .ce(N__47153),
            .sr(N__49361));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_10_6 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_10_6  (
            .in0(N__37241),
            .in1(N__41120),
            .in2(N__41319),
            .in3(N__37220),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_7 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_7  (
            .in0(N__32999),
            .in1(N__32982),
            .in2(N__32966),
            .in3(N__33354),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_11_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_11_1  (
            .in0(N__33293),
            .in1(N__33280),
            .in2(N__33263),
            .in3(N__33238),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_12_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_12_11_2  (
            .in0(N__33068),
            .in1(N__33027),
            .in2(_gnd_net_),
            .in3(N__36720),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49829),
            .ce(N__33334),
            .sr(N__49368));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_5 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_5  (
            .in0(N__32998),
            .in1(N__32981),
            .in2(N__32967),
            .in3(N__33353),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_12_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_12_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_12_11_6  (
            .in0(N__36230),
            .in1(N__36763),
            .in2(_gnd_net_),
            .in3(N__36719),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49829),
            .ce(N__33334),
            .sr(N__49368));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_12_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_12_0  (
            .in0(N__34383),
            .in1(N__35778),
            .in2(_gnd_net_),
            .in3(N__38490),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_12_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_12_12_1 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_12_12_1  (
            .in0(N__33294),
            .in1(N__33281),
            .in2(N__33264),
            .in3(N__33239),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_12_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_12_2  (
            .in0(N__34512),
            .in1(N__35754),
            .in2(_gnd_net_),
            .in3(N__38491),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_12_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_12_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_12_12_3  (
            .in0(N__33148),
            .in1(N__33202),
            .in2(_gnd_net_),
            .in3(N__36718),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_12_13_0  (
            .in0(N__46913),
            .in1(N__37901),
            .in2(_gnd_net_),
            .in3(N__39273),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49819),
            .ce(N__47152),
            .sr(N__49378));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_12_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_12_13_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_12_13_1  (
            .in0(N__39612),
            .in1(N__34345),
            .in2(_gnd_net_),
            .in3(N__46914),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49819),
            .ce(N__47152),
            .sr(N__49378));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_12_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_12_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_12_13_3  (
            .in0(N__39567),
            .in1(N__34453),
            .in2(_gnd_net_),
            .in3(N__46915),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49819),
            .ce(N__47152),
            .sr(N__49378));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_12_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_12_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_12_14_0  (
            .in0(N__34347),
            .in1(N__39611),
            .in2(_gnd_net_),
            .in3(N__46722),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_14_2 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_14_2  (
            .in0(N__34430),
            .in1(N__35478),
            .in2(N__35520),
            .in3(N__34416),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_12_14_3  (
            .in0(N__46723),
            .in1(N__37905),
            .in2(_gnd_net_),
            .in3(N__39272),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49817),
            .ce(N__37638),
            .sr(N__49382));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_15_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_15_0  (
            .in0(N__35910),
            .in1(N__34491),
            .in2(_gnd_net_),
            .in3(N__38460),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_15_1  (
            .in0(N__46830),
            .in1(N__34246),
            .in2(_gnd_net_),
            .in3(N__39653),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_15_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_15_2  (
            .in0(N__34455),
            .in1(N__39563),
            .in2(_gnd_net_),
            .in3(N__46831),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_15_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_15_3  (
            .in0(N__38462),
            .in1(N__35865),
            .in2(_gnd_net_),
            .in3(N__34626),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_15_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_15_4  (
            .in0(N__35850),
            .in1(N__34614),
            .in2(_gnd_net_),
            .in3(N__38463),
            .lcout(\current_shift_inst.control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_15_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_15_5  (
            .in0(N__38461),
            .in1(N__34470),
            .in2(_gnd_net_),
            .in3(N__35880),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_15_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_15_6  (
            .in0(N__34590),
            .in1(N__35826),
            .in2(_gnd_net_),
            .in3(N__38467),
            .lcout(\current_shift_inst.control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_15_7 .LUT_INIT=16'b0000010111110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_15_7  (
            .in0(N__34602),
            .in1(_gnd_net_),
            .in2(N__38492),
            .in3(N__35838),
            .lcout(\current_shift_inst.control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_12_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_12_16_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_12_16_0  (
            .in0(N__38493),
            .in1(N__35814),
            .in2(_gnd_net_),
            .in3(N__34578),
            .lcout(\current_shift_inst.control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_12_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_12_16_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_12_16_1  (
            .in0(N__38455),
            .in1(N__36000),
            .in2(_gnd_net_),
            .in3(N__34554),
            .lcout(\current_shift_inst.control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_16_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_16_2  (
            .in0(N__34542),
            .in1(N__35985),
            .in2(_gnd_net_),
            .in3(N__38456),
            .lcout(\current_shift_inst.control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_16_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_16_3  (
            .in0(N__38457),
            .in1(N__34530),
            .in2(_gnd_net_),
            .in3(N__35970),
            .lcout(\current_shift_inst.control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_16_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_16_4  (
            .in0(N__35895),
            .in1(N__34479),
            .in2(_gnd_net_),
            .in3(N__38454),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_16_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_16_6  (
            .in0(N__34695),
            .in1(N__35949),
            .in2(_gnd_net_),
            .in3(N__38458),
            .lcout(\current_shift_inst.control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_16_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_16_7  (
            .in0(N__38459),
            .in1(N__34683),
            .in2(_gnd_net_),
            .in3(N__35937),
            .lcout(\current_shift_inst.control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_1  (
            .in0(N__34671),
            .in1(N__35925),
            .in2(_gnd_net_),
            .in3(N__38494),
            .lcout(\current_shift_inst.control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2  (
            .in0(N__38495),
            .in1(N__34644),
            .in2(_gnd_net_),
            .in3(N__36078),
            .lcout(\current_shift_inst.control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_12_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_12_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_12_19_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_12_19_0  (
            .in0(N__49991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33543),
            .ce(),
            .sr(N__49404));
    defparam \delay_measurement_inst.start_timer_hc_LC_12_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49990),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33543),
            .ce(),
            .sr(N__49404));
    defparam \phase_controller_inst2.S1_LC_12_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_12_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33759),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49802),
            .ce(),
            .sr(N__49411));
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_0.C_ON=1'b0;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_0 (
            .in0(N__49476),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_red_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_13_2_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_13_2_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_13_2_1 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \phase_controller_inst1.state_3_LC_13_2_1  (
            .in0(N__35083),
            .in1(N__33452),
            .in2(N__33875),
            .in3(N__33504),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(),
            .sr(N__49291));
    defparam \phase_controller_inst1.state_2_LC_13_2_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_13_2_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_13_2_2 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.state_2_LC_13_2_2  (
            .in0(N__33809),
            .in1(N__33834),
            .in2(N__34910),
            .in3(N__33857),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(),
            .sr(N__49291));
    defparam \phase_controller_inst1.state_0_LC_13_2_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_13_2_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_13_2_3 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst1.state_0_LC_13_2_3  (
            .in0(N__34777),
            .in1(N__34727),
            .in2(N__33474),
            .in3(N__33497),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(),
            .sr(N__49291));
    defparam \phase_controller_inst1.state_4_LC_13_2_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_13_2_4 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_13_2_4 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_inst1.state_4_LC_13_2_4  (
            .in0(N__33453),
            .in1(N__33868),
            .in2(_gnd_net_),
            .in3(N__35084),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(),
            .sr(N__49291));
    defparam \phase_controller_inst1.start_flag_LC_13_2_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_flag_LC_13_2_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_flag_LC_13_2_5 .LUT_INIT=16'b1111100011111000;
    LogicCell40 \phase_controller_inst1.start_flag_LC_13_2_5  (
            .in0(N__35082),
            .in1(N__33451),
            .in2(N__33876),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.start_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(),
            .sr(N__49291));
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_13_3_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIE87F_2_LC_13_3_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \phase_controller_inst1.state_RNIE87F_2_LC_13_3_3  (
            .in0(N__33856),
            .in1(N__33828),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_3_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_3_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_3_5  (
            .in0(N__34778),
            .in1(N__33829),
            .in2(N__33858),
            .in3(N__34722),
            .lcout(\phase_controller_inst1.N_54_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36979),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49304));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_4_4 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_13_4_4  (
            .in0(N__33833),
            .in1(N__33948),
            .in2(N__37014),
            .in3(N__34142),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49304));
    defparam \phase_controller_inst1.start_timer_hc_LC_13_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_4_6 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_13_4_6  (
            .in0(N__33810),
            .in1(N__34745),
            .in2(N__34916),
            .in3(N__36978),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49304));
    defparam \phase_controller_inst2.state_3_LC_13_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_13_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_13_5_1 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \phase_controller_inst2.state_3_LC_13_5_1  (
            .in0(N__35087),
            .in1(N__35021),
            .in2(N__33768),
            .in3(N__35037),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49907),
            .ce(),
            .sr(N__49311));
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_13_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_13_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNIG7JF_2_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(N__38320),
            .in2(_gnd_net_),
            .in3(N__33725),
            .lcout(\phase_controller_inst2.N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_6_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__35718),
            .in2(_gnd_net_),
            .in3(N__35655),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_7_2 .LUT_INIT=16'b1011001110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_13_7_2  (
            .in0(N__33960),
            .in1(N__37012),
            .in2(N__34143),
            .in3(N__33944),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49882),
            .ce(),
            .sr(N__49326));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_13_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_13_7_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_13_7_3  (
            .in0(N__37011),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34138),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33963),
            .in3(N__33942),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_7_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_7_5  (
            .in0(N__37010),
            .in1(N__33959),
            .in2(_gnd_net_),
            .in3(N__36980),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_13_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_13_7_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33951),
            .in3(N__33923),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_7_7 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_7_7  (
            .in0(N__33943),
            .in1(N__37590),
            .in2(N__33927),
            .in3(N__34946),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49882),
            .ce(),
            .sr(N__49326));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_13_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_13_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__37107),
            .in2(N__33915),
            .in3(N__34942),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_13_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_13_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__37095),
            .in2(N__33906),
            .in3(N__35234),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_13_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_13_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_13_8_2  (
            .in0(N__35210),
            .in1(N__34365),
            .in2(N__33897),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_13_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_13_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__37659),
            .in2(N__33885),
            .in3(N__35195),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_13_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_13_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__34974),
            .in2(N__34050),
            .in3(N__35180),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_13_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_13_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__34038),
            .in2(N__34098),
            .in3(N__35165),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_13_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_13_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__34191),
            .in2(N__34032),
            .in3(N__35150),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_13_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_13_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__34023),
            .in2(N__34011),
            .in3(N__35135),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_13_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_13_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__34170),
            .in2(N__33999),
            .in3(N__35120),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_13_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_13_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__33990),
            .in2(N__34311),
            .in3(N__35333),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_13_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_13_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_13_9_2  (
            .in0(N__35318),
            .in1(N__34329),
            .in2(N__33984),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_13_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_13_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_13_9_3  (
            .in0(N__35303),
            .in1(N__34356),
            .in2(N__33972),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_13_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_13_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__34074),
            .in2(N__35424),
            .in3(N__35288),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_13_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_13_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__36939),
            .in2(N__34068),
            .in3(N__35273),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_13_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_13_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__34182),
            .in2(N__34059),
            .in3(N__35258),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_13_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_13_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__36864),
            .in2(N__36927),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_13_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_13_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__37284),
            .in2(N__37083),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_13_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_13_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__37146),
            .in2(N__37029),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_13_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_13_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__37716),
            .in2(N__37776),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_13_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_13_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__34989),
            .in2(N__35004),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_13_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_13_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__34107),
            .in2(N__34116),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_13_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_13_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__34200),
            .in2(N__34281),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_13_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_13_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__34158),
            .in2(N__34404),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_13_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_13_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34146),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_13_11_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_13_11_0  (
            .in0(N__35351),
            .in1(N__34290),
            .in2(N__34086),
            .in3(N__35581),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_13_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_13_11_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_13_11_1  (
            .in0(N__34289),
            .in1(N__34085),
            .in2(N__35583),
            .in3(N__35350),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_13_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_13_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_13_11_3  (
            .in0(N__46849),
            .in1(N__45443),
            .in2(_gnd_net_),
            .in3(N__45407),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(elapsed_time_ns_1_RNII43T9_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_13_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_13_11_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_13_11_4  (
            .in0(N__45444),
            .in1(_gnd_net_),
            .in2(N__34101),
            .in3(N__46853),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(N__37607),
            .sr(N__49362));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_13_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_13_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_13_11_5  (
            .in0(N__46852),
            .in1(N__47121),
            .in2(_gnd_net_),
            .in3(N__50382),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(N__37607),
            .sr(N__49362));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_11_6  (
            .in0(N__41630),
            .in1(N__41597),
            .in2(_gnd_net_),
            .in3(N__46850),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(elapsed_time_ns_1_RNI47DN9_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_13_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_13_11_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_13_11_7  (
            .in0(N__46851),
            .in1(_gnd_net_),
            .in2(N__34293),
            .in3(N__41631),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(N__37607),
            .sr(N__49362));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_12_0 .LUT_INIT=16'b0111001100010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_12_0  (
            .in0(N__35562),
            .in1(N__35541),
            .in2(N__34224),
            .in3(N__34209),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_12_1  (
            .in0(N__46814),
            .in1(N__39694),
            .in2(_gnd_net_),
            .in3(N__34265),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(elapsed_time_ns_1_RNI69DN9_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_13_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_13_12_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_13_12_2  (
            .in0(N__39695),
            .in1(_gnd_net_),
            .in2(N__34254),
            .in3(N__46816),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49831),
            .ce(N__37608),
            .sr(N__49369));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_13_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_13_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_13_12_3  (
            .in0(N__46815),
            .in1(N__34251),
            .in2(_gnd_net_),
            .in3(N__39649),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49831),
            .ce(N__37608),
            .sr(N__49369));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_12_4 .LUT_INIT=16'b1111011100110001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_12_4  (
            .in0(N__35561),
            .in1(N__35540),
            .in2(N__34223),
            .in3(N__34208),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_13_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_13_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_13_12_6  (
            .in0(N__45383),
            .in1(N__45354),
            .in2(_gnd_net_),
            .in3(N__46817),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49831),
            .ce(N__37608),
            .sr(N__49369));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_13_13_0  (
            .in0(N__46916),
            .in1(N__45208),
            .in2(_gnd_net_),
            .in3(N__45191),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(N__37641),
            .sr(N__49373));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_13_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_13_13_1  (
            .in0(N__41400),
            .in1(N__46921),
            .in2(_gnd_net_),
            .in3(N__41433),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(N__37641),
            .sr(N__49373));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_13_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_13_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_13_13_2  (
            .in0(N__46918),
            .in1(N__41475),
            .in2(_gnd_net_),
            .in3(N__41514),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(N__37641),
            .sr(N__49373));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_3  (
            .in0(N__41343),
            .in1(N__46920),
            .in2(_gnd_net_),
            .in3(N__41376),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(N__37641),
            .sr(N__49373));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_13_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_13_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_13_13_4  (
            .in0(N__46917),
            .in1(N__39600),
            .in2(_gnd_net_),
            .in3(N__34346),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(N__37641),
            .sr(N__49373));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_13_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_13_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_13_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_13_13_5  (
            .in0(N__40921),
            .in1(N__46919),
            .in2(_gnd_net_),
            .in3(N__40961),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(N__37641),
            .sr(N__49373));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_14_0  (
            .in0(N__41375),
            .in1(N__40996),
            .in2(N__40962),
            .in3(N__41432),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_14_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_14_1  (
            .in0(N__45442),
            .in1(N__39316),
            .in2(N__34320),
            .in3(N__34317),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_14_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__39268),
            .in2(_gnd_net_),
            .in3(N__45353),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_13_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_13_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_13_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_13_14_3  (
            .in0(N__40997),
            .in1(N__41024),
            .in2(_gnd_net_),
            .in3(N__46724),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49820),
            .ce(N__37639),
            .sr(N__49379));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_15_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_15_5  (
            .in0(N__35439),
            .in1(N__34299),
            .in2(N__35733),
            .in3(N__39561),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_13_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_13_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_13_15_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_13_15_6  (
            .in0(N__39562),
            .in1(_gnd_net_),
            .in2(N__34458),
            .in3(N__34454),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49818),
            .ce(N__37642),
            .sr(N__49383));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_13_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_13_15_7 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_13_15_7  (
            .in0(N__34431),
            .in1(N__35477),
            .in2(N__35519),
            .in3(N__34415),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_13_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_13_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__36795),
            .in2(N__41883),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_13_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_13_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__46369),
            .in2(N__46338),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_13_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_13_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__47641),
            .in2(N__37959),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_13_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_13_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__39504),
            .in2(N__47807),
            .in3(N__34389),
            .lcout(\current_shift_inst.un38_control_input_0_s1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_13_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_13_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(N__47645),
            .in2(N__39777),
            .in3(N__34386),
            .lcout(\current_shift_inst.un38_control_input_0_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_13_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_13_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(N__39897),
            .in2(N__47808),
            .in3(N__34371),
            .lcout(\current_shift_inst.un38_control_input_0_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_13_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_13_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__47649),
            .in2(N__38133),
            .in3(N__34368),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_13_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_13_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(N__36039),
            .in2(N__47809),
            .in3(N__34518),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_13_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_13_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__47653),
            .in2(N__36171),
            .in3(N__34515),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_13_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_13_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__39738),
            .in2(N__47810),
            .in3(N__34500),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_13_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_13_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__47657),
            .in2(N__48336),
            .in3(N__34497),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_13_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_13_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__36162),
            .in2(N__47811),
            .in3(N__34494),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_13_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_13_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__47661),
            .in2(N__48405),
            .in3(N__34482),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_13_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_13_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__47253),
            .in2(N__47812),
            .in3(N__34473),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_13_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_13_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__47665),
            .in2(N__38217),
            .in3(N__34461),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_13_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_13_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__39789),
            .in2(N__47813),
            .in3(N__34617),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_13_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_13_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__47685),
            .in2(N__36834),
            .in3(N__34605),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_13_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__36024),
            .in2(N__47818),
            .in3(N__34593),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_13_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_13_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__47689),
            .in2(N__36033),
            .in3(N__34581),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_13_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_13_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__36012),
            .in2(N__47819),
            .in3(N__34569),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_13_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_13_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__47693),
            .in2(N__39939),
            .in3(N__34557),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_13_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_13_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__36018),
            .in2(N__47820),
            .in3(N__34545),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_13_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_13_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__47697),
            .in2(N__39966),
            .in3(N__34533),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_13_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_13_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__36147),
            .in2(N__47821),
            .in3(N__34521),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_13_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_13_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__47822),
            .in2(N__36843),
            .in3(N__34701),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_13_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_13_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__42621),
            .in2(N__47872),
            .in3(N__34698),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_13_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_13_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__47826),
            .in2(N__36852),
            .in3(N__34686),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_13_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_13_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__36132),
            .in2(N__47873),
            .in3(N__34674),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_13_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_13_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__47830),
            .in2(N__36156),
            .in3(N__34662),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_13_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_13_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__36126),
            .in2(N__47874),
            .in3(N__34647),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_13_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_13_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__47834),
            .in2(N__36141),
            .in3(N__34632),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_13_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_13_19_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_13_19_7  (
            .in0(N__47835),
            .in1(N__48255),
            .in2(_gnd_net_),
            .in3(N__34629),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34734),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(N__49412));
    defparam \current_shift_inst.start_timer_s1_LC_13_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_13_22_4 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_22_4  (
            .in0(N__34855),
            .in1(N__34836),
            .in2(_gnd_net_),
            .in3(N__34914),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(N__49412));
    defparam \phase_controller_inst1.S1_LC_13_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34915),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(N__49412));
    defparam \current_shift_inst.stop_timer_s1_LC_13_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_13_23_4 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_23_4  (
            .in0(N__34837),
            .in1(N__34815),
            .in2(N__34917),
            .in3(N__34856),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49800),
            .ce(),
            .sr(N__49417));
    defparam \current_shift_inst.timer_s1.running_LC_13_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_23_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_23_7  (
            .in0(N__34814),
            .in1(N__34838),
            .in2(_gnd_net_),
            .in3(N__36198),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49800),
            .ce(),
            .sr(N__49417));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_24_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_24_4  (
            .in0(N__36196),
            .in1(N__34813),
            .in2(_gnd_net_),
            .in3(N__34839),
            .lcout(\current_shift_inst.timer_s1.N_162_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__36195),
            .in2(_gnd_net_),
            .in3(N__34812),
            .lcout(\current_shift_inst.timer_s1.N_161_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_14_3_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_14_3_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_14_3_0 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \phase_controller_inst1.state_1_LC_14_3_0  (
            .in0(N__34782),
            .in1(N__34746),
            .in2(_gnd_net_),
            .in3(N__34726),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49941),
            .ce(),
            .sr(N__49292));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_14_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_14_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_14_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38984),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49930),
            .ce(),
            .sr(N__49296));
    defparam \phase_controller_inst2.state_4_LC_14_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_4_LC_14_5_1 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst2.state_4_LC_14_5_1 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_inst2.state_4_LC_14_5_1  (
            .in0(N__35035),
            .in1(N__35017),
            .in2(_gnd_net_),
            .in3(N__35086),
            .lcout(\phase_controller_inst2.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49919),
            .ce(),
            .sr(N__49305));
    defparam \phase_controller_inst2.start_flag_LC_14_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_flag_LC_14_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_flag_LC_14_5_2 .LUT_INIT=16'b1111100011111000;
    LogicCell40 \phase_controller_inst2.start_flag_LC_14_5_2  (
            .in0(N__35085),
            .in1(N__35036),
            .in2(N__35022),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.start_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49919),
            .ce(),
            .sr(N__49305));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_6_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_6_0  (
            .in0(N__35396),
            .in1(N__34962),
            .in2(N__36954),
            .in3(N__35375),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_6_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_6_1  (
            .in0(N__34961),
            .in1(N__35397),
            .in2(N__35376),
            .in3(N__36953),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_14_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_14_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_14_6_2  (
            .in0(N__45038),
            .in1(N__45014),
            .in2(_gnd_net_),
            .in3(N__46956),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_3  (
            .in0(N__46957),
            .in1(N__39317),
            .in2(_gnd_net_),
            .in3(N__37040),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(elapsed_time_ns_1_RNIH33T9_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_14_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_14_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_14_6_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_14_6_4  (
            .in0(N__39318),
            .in1(_gnd_net_),
            .in2(N__34977),
            .in3(N__46960),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49908),
            .ce(N__37643),
            .sr(N__49312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_6_6  (
            .in0(N__40477),
            .in1(N__46958),
            .in2(_gnd_net_),
            .in3(N__40436),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(elapsed_time_ns_1_RNI25DN9_0_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_14_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_14_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_14_6_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_14_6_7  (
            .in0(N__46959),
            .in1(_gnd_net_),
            .in2(N__34965),
            .in3(N__40478),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49908),
            .ce(N__37643),
            .sr(N__49312));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__34953),
            .in2(N__34947),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_7_1  (
            .in0(N__37506),
            .in1(N__35235),
            .in2(_gnd_net_),
            .in3(N__35223),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_7_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_7_2  (
            .in0(N__37587),
            .in1(N__35211),
            .in2(N__35220),
            .in3(N__35199),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_14_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_14_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_14_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_14_7_3  (
            .in0(N__37507),
            .in1(N__35196),
            .in2(_gnd_net_),
            .in3(N__35184),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_14_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_14_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_14_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_14_7_4  (
            .in0(N__37588),
            .in1(N__35181),
            .in2(_gnd_net_),
            .in3(N__35169),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_7_5  (
            .in0(N__37508),
            .in1(N__35166),
            .in2(_gnd_net_),
            .in3(N__35154),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_14_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_14_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_14_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_14_7_6  (
            .in0(N__37589),
            .in1(N__35151),
            .in2(_gnd_net_),
            .in3(N__35139),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_7_7  (
            .in0(N__37509),
            .in1(N__35136),
            .in2(_gnd_net_),
            .in3(N__35124),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49897),
            .ce(),
            .sr(N__49319));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_14_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_14_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_14_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_14_8_0  (
            .in0(N__37586),
            .in1(N__35121),
            .in2(_gnd_net_),
            .in3(N__35109),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49883),
            .ce(),
            .sr(N__49327));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_8_1  (
            .in0(N__37555),
            .in1(N__35334),
            .in2(_gnd_net_),
            .in3(N__35322),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49883),
            .ce(),
            .sr(N__49327));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_8_2  (
            .in0(N__37583),
            .in1(N__35319),
            .in2(_gnd_net_),
            .in3(N__35307),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49883),
            .ce(),
            .sr(N__49327));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_8_3  (
            .in0(N__37556),
            .in1(N__35304),
            .in2(_gnd_net_),
            .in3(N__35292),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49883),
            .ce(),
            .sr(N__49327));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_14_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_14_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_14_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_14_8_4  (
            .in0(N__37584),
            .in1(N__35289),
            .in2(_gnd_net_),
            .in3(N__35277),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49883),
            .ce(),
            .sr(N__49327));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_8_5  (
            .in0(N__37557),
            .in1(N__35274),
            .in2(_gnd_net_),
            .in3(N__35262),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49883),
            .ce(),
            .sr(N__49327));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_8_6  (
            .in0(N__37585),
            .in1(N__35259),
            .in2(_gnd_net_),
            .in3(N__35247),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49883),
            .ce(),
            .sr(N__49327));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_8_7  (
            .in0(N__37558),
            .in1(N__36912),
            .in2(_gnd_net_),
            .in3(N__35244),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49883),
            .ce(),
            .sr(N__49327));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_9_0  (
            .in0(N__37622),
            .in1(N__36880),
            .in2(_gnd_net_),
            .in3(N__35241),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49873),
            .ce(),
            .sr(N__49335));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_9_1  (
            .in0(N__37609),
            .in1(N__37299),
            .in2(_gnd_net_),
            .in3(N__35238),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49873),
            .ce(),
            .sr(N__49335));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_14_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_14_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_14_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_14_9_2  (
            .in0(N__37623),
            .in1(N__37329),
            .in2(_gnd_net_),
            .in3(N__35412),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49873),
            .ce(),
            .sr(N__49335));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_14_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_14_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_14_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_14_9_3  (
            .in0(N__37610),
            .in1(N__37163),
            .in2(_gnd_net_),
            .in3(N__35409),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49873),
            .ce(),
            .sr(N__49335));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_14_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_14_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_14_9_4  (
            .in0(N__37624),
            .in1(N__37179),
            .in2(_gnd_net_),
            .in3(N__35406),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49873),
            .ce(),
            .sr(N__49335));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_14_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_14_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_14_9_5  (
            .in0(N__37611),
            .in1(N__37753),
            .in2(_gnd_net_),
            .in3(N__35403),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49873),
            .ce(),
            .sr(N__49335));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_14_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_14_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_14_9_6  (
            .in0(N__37625),
            .in1(N__37732),
            .in2(_gnd_net_),
            .in3(N__35400),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49873),
            .ce(),
            .sr(N__49335));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_14_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_14_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_14_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_14_9_7  (
            .in0(N__37612),
            .in1(N__35395),
            .in2(_gnd_net_),
            .in3(N__35379),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49873),
            .ce(),
            .sr(N__49335));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_14_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_14_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_14_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_14_10_0  (
            .in0(N__37619),
            .in1(N__35371),
            .in2(_gnd_net_),
            .in3(N__35355),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49345));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_14_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_14_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_14_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_14_10_1  (
            .in0(N__37626),
            .in1(N__35352),
            .in2(_gnd_net_),
            .in3(N__35337),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49345));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_14_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_14_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_14_10_2  (
            .in0(N__37620),
            .in1(N__35582),
            .in2(_gnd_net_),
            .in3(N__35565),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49345));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_14_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_14_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_14_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_14_10_3  (
            .in0(N__37627),
            .in1(N__35560),
            .in2(_gnd_net_),
            .in3(N__35544),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49345));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_14_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_14_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_14_10_4  (
            .in0(N__37621),
            .in1(N__35539),
            .in2(_gnd_net_),
            .in3(N__35523),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49345));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_14_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_14_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_14_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_14_10_5  (
            .in0(N__37628),
            .in1(N__35506),
            .in2(_gnd_net_),
            .in3(N__35484),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49345));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_14_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_14_10_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_14_10_6  (
            .in0(N__35470),
            .in1(N__37629),
            .in2(_gnd_net_),
            .in3(N__35481),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49863),
            .ce(),
            .sr(N__49345));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_14_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_14_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_14_11_2  (
            .in0(N__39464),
            .in1(N__44663),
            .in2(N__47243),
            .in3(N__44574),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_14_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_14_11_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_14_11_3  (
            .in0(N__41558),
            .in1(N__41682),
            .in2(N__45516),
            .in3(N__40468),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_14_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_14_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_14_11_4  (
            .in0(N__35589),
            .in1(N__35448),
            .in2(N__35442),
            .in3(N__37269),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_14_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_14_11_6  (
            .in0(N__44354),
            .in1(N__44321),
            .in2(_gnd_net_),
            .in3(N__46936),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49851),
            .ce(N__37630),
            .sr(N__49354));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_12_0  (
            .in0(N__46812),
            .in1(N__37679),
            .in2(_gnd_net_),
            .in3(N__39353),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_14_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_14_12_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_14_12_1  (
            .in0(N__39693),
            .in1(N__37275),
            .in2(_gnd_net_),
            .in3(N__47112),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_12_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_12_4  (
            .in0(N__46813),
            .in1(N__40925),
            .in2(_gnd_net_),
            .in3(N__40960),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_12_5  (
            .in0(N__45212),
            .in1(N__45190),
            .in2(_gnd_net_),
            .in3(N__46811),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_12_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_12_6  (
            .in0(N__35717),
            .in1(N__35679),
            .in2(_gnd_net_),
            .in3(N__35661),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_12_7  (
            .in0(N__39648),
            .in1(N__41624),
            .in2(N__39610),
            .in3(N__45003),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__36794),
            .in2(N__41445),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__46359),
            .in2(N__41853),
            .in3(N__38271),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2  (
            .in0(N__38272),
            .in1(N__47379),
            .in2(N__37380),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__37815),
            .in2(N__47584),
            .in3(N__35784),
            .lcout(\current_shift_inst.un38_control_input_0_s0_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__47383),
            .in2(N__41802),
            .in3(N__35781),
            .lcout(\current_shift_inst.un38_control_input_0_s0_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__39750),
            .in2(N__47585),
            .in3(N__35766),
            .lcout(\current_shift_inst.un38_control_input_0_s0_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__47387),
            .in2(N__37983),
            .in3(N__35763),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__37800),
            .in2(N__47586),
            .in3(N__35760),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__47391),
            .in2(N__37932),
            .in3(N__35757),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__37923),
            .in2(N__47587),
            .in3(N__35742),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__47395),
            .in2(N__37809),
            .in3(N__35739),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__37785),
            .in2(N__47588),
            .in3(N__35736),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__47399),
            .in2(N__37794),
            .in3(N__35898),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__39909),
            .in2(N__47589),
            .in3(N__35883),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__47403),
            .in2(N__37974),
            .in3(N__35868),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__37965),
            .in2(N__47590),
            .in3(N__35853),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__47669),
            .in2(N__38088),
            .in3(N__35841),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__37917),
            .in2(N__47814),
            .in3(N__35829),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__47673),
            .in2(N__38010),
            .in3(N__35817),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__37911),
            .in2(N__47815),
            .in3(N__35802),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__47677),
            .in2(N__48270),
            .in3(N__35787),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__38205),
            .in2(N__47816),
            .in3(N__35988),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__47681),
            .in2(N__37944),
            .in3(N__35973),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__38226),
            .in2(N__47817),
            .in3(N__35958),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__36006),
            .in2(N__47836),
            .in3(N__35955),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__47721),
            .in2(N__38196),
            .in3(N__35952),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__37992),
            .in2(N__47837),
            .in3(N__35940),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__47725),
            .in2(N__38187),
            .in3(N__35928),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__36177),
            .in2(N__47838),
            .in3(N__35913),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__47729),
            .in2(N__38175),
            .in3(N__36081),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__37998),
            .in2(N__47839),
            .in3(N__36066),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7  (
            .in0(N__46590),
            .in1(N__36063),
            .in2(N__38499),
            .in3(N__36051),
            .lcout(\current_shift_inst.control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_14_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_14_17_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_14_17_0  (
            .in0(N__48208),
            .in1(N__47741),
            .in2(N__40037),
            .in3(N__42009),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_14_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_14_17_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_14_17_1  (
            .in0(N__47739),
            .in1(N__48211),
            .in2(N__42180),
            .in3(N__43164),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_14_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_14_17_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_14_17_2  (
            .in0(N__48210),
            .in1(N__47746),
            .in2(N__40562),
            .in3(N__42211),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_14_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_14_17_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_14_17_3  (
            .in0(N__47743),
            .in1(N__48213),
            .in2(N__42093),
            .in3(N__40326),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_14_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_14_17_4 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_14_17_4  (
            .in0(N__48212),
            .in1(N__42140),
            .in2(N__42612),
            .in3(N__47744),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_17_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_17_5  (
            .in0(N__47745),
            .in1(N__48214),
            .in2(N__43061),
            .in3(N__42485),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_17_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_17_6  (
            .in0(N__48215),
            .in1(N__47740),
            .in2(N__43014),
            .in3(N__42389),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_14_17_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_14_17_7  (
            .in0(N__47742),
            .in1(N__48209),
            .in2(N__42713),
            .in3(N__41976),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_14_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_14_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_14_18_0  (
            .in0(N__48216),
            .in1(N__43382),
            .in2(N__47847),
            .in3(N__43344),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_18_1 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_18_1  (
            .in0(N__42390),
            .in1(N__47750),
            .in2(N__43013),
            .in3(N__48222),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_14_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_14_18_2 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_14_18_2  (
            .in0(N__47754),
            .in1(N__42519),
            .in2(N__48251),
            .in3(N__40221),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_14_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_14_18_3 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_14_18_3  (
            .in0(N__42310),
            .in1(N__47757),
            .in2(N__38277),
            .in3(N__48224),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_4  (
            .in0(N__48221),
            .in1(N__42419),
            .in2(N__47846),
            .in3(N__42908),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_14_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_14_18_5 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_14_18_5  (
            .in0(N__42353),
            .in1(N__47755),
            .in2(N__43532),
            .in3(N__48223),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_18_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_18_6  (
            .in0(N__36120),
            .in1(N__36111),
            .in2(_gnd_net_),
            .in3(N__38485),
            .lcout(\current_shift_inst.control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_7 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_7  (
            .in0(N__42457),
            .in1(N__47756),
            .in2(N__42959),
            .in3(N__48220),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_14_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_14_19_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_14_19_1  (
            .in0(N__47870),
            .in1(N__48253),
            .in2(N__43062),
            .in3(N__42489),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_14_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_14_19_2 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_14_19_2  (
            .in0(N__48252),
            .in1(N__42249),
            .in2(N__43260),
            .in3(N__47871),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3  (
            .in0(N__38442),
            .in1(N__36822),
            .in2(_gnd_net_),
            .in3(N__36816),
            .lcout(\current_shift_inst.control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_20_0  (
            .in0(N__41882),
            .in1(N__38754),
            .in2(_gnd_net_),
            .in3(N__38253),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_14_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_14_20_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_14_20_3  (
            .in0(N__36223),
            .in1(N__36774),
            .in2(_gnd_net_),
            .in3(N__36723),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_21_2  (
            .in0(N__46553),
            .in1(N__38753),
            .in2(_gnd_net_),
            .in3(N__36204),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_21_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__46525),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49809),
            .ce(N__46406),
            .sr(N__49405));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36197),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_15_4_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_15_4_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_15_4_1  (
            .in0(N__39001),
            .in1(N__38291),
            .in2(_gnd_net_),
            .in3(N__38980),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_15_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_15_4_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__37013),
            .in2(_gnd_net_),
            .in3(N__36981),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_15_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_15_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_15_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_15_5_3  (
            .in0(N__44589),
            .in1(N__44612),
            .in2(_gnd_net_),
            .in3(N__47038),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49931),
            .ce(N__37518),
            .sr(N__49297));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_15_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_15_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_15_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_15_6_1  (
            .in0(N__45034),
            .in1(N__47076),
            .in2(_gnd_net_),
            .in3(N__45015),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49920),
            .ce(N__37644),
            .sr(N__49306));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0  (
            .in0(N__44545),
            .in1(N__44513),
            .in2(_gnd_net_),
            .in3(N__47029),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(elapsed_time_ns_1_RNI13CN9_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_15_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_15_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_15_7_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_15_7_1  (
            .in0(N__47030),
            .in1(_gnd_net_),
            .in2(N__36942),
            .in3(N__44546),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49909),
            .ce(N__37597),
            .sr(N__49313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_15_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_15_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_15_7_2  (
            .in0(N__44611),
            .in1(N__44584),
            .in2(_gnd_net_),
            .in3(N__47028),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_15_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_15_7_4 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_15_7_4  (
            .in0(N__36881),
            .in1(N__37067),
            .in2(N__36897),
            .in3(N__36910),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_7_5 .LUT_INIT=16'b0100000011011100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_7_5  (
            .in0(N__36911),
            .in1(N__36893),
            .in2(N__37068),
            .in3(N__36882),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_15_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_15_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_15_7_6  (
            .in0(N__44416),
            .in1(N__47027),
            .in2(_gnd_net_),
            .in3(N__44375),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(elapsed_time_ns_1_RNI35CN9_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_15_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_15_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_15_7_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_15_7_7  (
            .in0(N__47031),
            .in1(_gnd_net_),
            .in2(N__37071),
            .in3(N__44417),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49909),
            .ce(N__37597),
            .sr(N__49313));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_8_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_8_0  (
            .in0(N__40710),
            .in1(N__40733),
            .in2(N__37056),
            .in3(N__47190),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_8_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_8_1  (
            .in0(N__47189),
            .in1(N__40709),
            .in2(N__40737),
            .in3(N__37052),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_15_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_15_8_3  (
            .in0(N__37263),
            .in1(N__39465),
            .in2(_gnd_net_),
            .in3(N__47035),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49898),
            .ce(N__47156),
            .sr(N__49320));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_15_8_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_15_8_4  (
            .in0(N__47033),
            .in1(N__37200),
            .in2(N__39537),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49898),
            .ce(N__47156),
            .sr(N__49320));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_15_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_15_8_5  (
            .in0(N__41474),
            .in1(N__41509),
            .in2(_gnd_net_),
            .in3(N__47036),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49898),
            .ce(N__47156),
            .sr(N__49320));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_15_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_15_8_6  (
            .in0(N__47034),
            .in1(N__37683),
            .in2(_gnd_net_),
            .in3(N__39352),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49898),
            .ce(N__47156),
            .sr(N__49320));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_15_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_15_8_7  (
            .in0(N__37044),
            .in1(N__39315),
            .in2(_gnd_net_),
            .in3(N__47037),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49898),
            .ce(N__47156),
            .sr(N__49320));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_9_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_9_0  (
            .in0(N__37178),
            .in1(N__37159),
            .in2(N__37131),
            .in3(N__37116),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_15_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_15_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_15_9_1  (
            .in0(N__37115),
            .in1(N__37177),
            .in2(N__37164),
            .in3(N__37130),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_15_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_15_9_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_15_9_2  (
            .in0(N__46965),
            .in1(_gnd_net_),
            .in2(N__45514),
            .in3(N__45467),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(elapsed_time_ns_1_RNIV1DN9_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_15_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_15_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_15_9_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__45507),
            .in2(N__37134),
            .in3(N__46970),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49884),
            .ce(N__37519),
            .sr(N__49328));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_9_4  (
            .in0(N__46964),
            .in1(N__44661),
            .in2(_gnd_net_),
            .in3(N__44624),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_15_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_15_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_15_9_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_15_9_5  (
            .in0(N__44662),
            .in1(_gnd_net_),
            .in2(N__37119),
            .in3(N__46969),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49884),
            .ce(N__37519),
            .sr(N__49328));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_15_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_15_9_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_15_9_6  (
            .in0(N__50325),
            .in1(_gnd_net_),
            .in2(N__47039),
            .in3(N__45146),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49884),
            .ce(N__37519),
            .sr(N__49328));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_15_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_15_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_15_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_15_9_7  (
            .in0(N__37199),
            .in1(N__39533),
            .in2(_gnd_net_),
            .in3(N__46971),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49884),
            .ce(N__37519),
            .sr(N__49328));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_10_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_10_0  (
            .in0(N__37338),
            .in1(N__37328),
            .in2(N__37313),
            .in3(N__37298),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_10_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_10_1  (
            .in0(N__47232),
            .in1(N__47058),
            .in2(_gnd_net_),
            .in3(N__47201),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(elapsed_time_ns_1_RNI57CN9_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_15_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_15_10_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_15_10_2  (
            .in0(N__47059),
            .in1(_gnd_net_),
            .in2(N__37341),
            .in3(N__47233),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49874),
            .ce(N__37634),
            .sr(N__49336));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_15_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_15_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_15_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_15_10_3  (
            .in0(N__37258),
            .in1(N__39460),
            .in2(_gnd_net_),
            .in3(N__47060),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49874),
            .ce(N__37634),
            .sr(N__49336));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_15_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_15_10_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_15_10_4  (
            .in0(N__37337),
            .in1(N__37327),
            .in2(N__37314),
            .in3(N__37297),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_11_0  (
            .in0(N__41496),
            .in1(N__39337),
            .in2(N__39532),
            .in3(N__50319),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_11_1  (
            .in0(N__45172),
            .in1(N__44530),
            .in2(N__44407),
            .in3(N__44310),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_11_2  (
            .in0(N__37262),
            .in1(N__39450),
            .in2(_gnd_net_),
            .in3(N__46934),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_11_4 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_11_4  (
            .in0(N__37242),
            .in1(N__41318),
            .in2(N__41127),
            .in3(N__37221),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_5  (
            .in0(N__46935),
            .in1(N__37198),
            .in2(_gnd_net_),
            .in3(N__39525),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_15_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_15_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_15_11_7  (
            .in0(N__46933),
            .in1(N__45376),
            .in2(_gnd_net_),
            .in3(N__45342),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_15_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_15_12_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_15_12_0  (
            .in0(N__37704),
            .in1(N__37692),
            .in2(N__37758),
            .in3(N__37736),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_15_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_15_12_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_15_12_1  (
            .in0(N__37691),
            .in1(N__37757),
            .in2(N__37737),
            .in3(N__37703),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_15_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_15_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_15_12_3  (
            .in0(N__46942),
            .in1(N__41585),
            .in2(_gnd_net_),
            .in3(N__41550),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49852),
            .ce(N__37640),
            .sr(N__49355));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_15_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_15_12_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_15_12_4  (
            .in0(N__41676),
            .in1(N__46940),
            .in2(_gnd_net_),
            .in3(N__41651),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(elapsed_time_ns_1_RNI03DN9_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_15_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_15_12_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_15_12_5  (
            .in0(N__46941),
            .in1(_gnd_net_),
            .in2(N__37695),
            .in3(N__41677),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49852),
            .ce(N__37640),
            .sr(N__49355));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_15_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_15_12_7  (
            .in0(N__46943),
            .in1(N__37675),
            .in2(_gnd_net_),
            .in3(N__39354),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49852),
            .ce(N__37640),
            .sr(N__49355));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_13_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_13_0  (
            .in0(N__48093),
            .in1(N__47419),
            .in2(N__40095),
            .in3(N__41778),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_13_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_13_3  (
            .in0(N__38427),
            .in1(N__37371),
            .in2(_gnd_net_),
            .in3(N__37365),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_13_4  (
            .in0(N__39264),
            .in1(N__37900),
            .in2(_gnd_net_),
            .in3(N__46881),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_13_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_13_5  (
            .in0(N__38428),
            .in1(N__37881),
            .in2(_gnd_net_),
            .in3(N__37866),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_15_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_15_13_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_15_13_6  (
            .in0(N__37848),
            .in1(N__37842),
            .in2(_gnd_net_),
            .in3(N__38426),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_15_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_15_13_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_15_13_7  (
            .in0(N__47418),
            .in1(N__48094),
            .in2(N__42870),
            .in3(N__41751),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_14_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_14_0  (
            .in0(N__48393),
            .in1(N__48166),
            .in2(N__47610),
            .in3(N__48360),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_15_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_15_14_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_15_14_1  (
            .in0(N__48165),
            .in1(N__47426),
            .in2(N__40041),
            .in3(N__42008),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_14_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_14_2  (
            .in0(N__47428),
            .in1(N__48168),
            .in2(N__48432),
            .in3(N__48467),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_14_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_14_3  (
            .in0(N__41023),
            .in1(N__41001),
            .in2(_gnd_net_),
            .in3(N__46912),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_14_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_14_4  (
            .in0(N__47427),
            .in1(N__48167),
            .in2(N__43383),
            .in3(N__43343),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_14_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_14_6  (
            .in0(N__42759),
            .in1(N__48164),
            .in2(N__47611),
            .in3(N__42053),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_14_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_14_7  (
            .in0(N__48169),
            .in1(N__47429),
            .in2(N__43448),
            .in3(N__43485),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_15_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_15_15_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_15_15_1  (
            .in0(N__47616),
            .in1(N__48082),
            .in2(N__43110),
            .in3(N__42279),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_15_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_15_2  (
            .in0(N__48079),
            .in1(N__47618),
            .in2(N__40094),
            .in3(N__41774),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_15_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_15_3  (
            .in0(N__47614),
            .in1(N__48085),
            .in2(N__40263),
            .in3(N__42558),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_15_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_15_15_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_15_15_4  (
            .in0(N__48080),
            .in1(N__47613),
            .in2(N__42714),
            .in3(N__41972),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_15_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_15_15_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_15_15_5  (
            .in0(N__47612),
            .in1(N__48081),
            .in2(N__40170),
            .in3(N__41943),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_15_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_15_15_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_15_15_6  (
            .in0(N__48083),
            .in1(N__47617),
            .in2(N__40563),
            .in3(N__42213),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_15_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_15_7  (
            .in0(N__47615),
            .in1(N__48084),
            .in2(N__42141),
            .in3(N__42605),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_16_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_16_0  (
            .in0(N__38163),
            .in1(N__38154),
            .in2(_gnd_net_),
            .in3(N__38430),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_15_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_15_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_15_16_1  (
            .in0(N__48207),
            .in1(N__42758),
            .in2(N__47795),
            .in3(N__42054),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_16_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_16_2  (
            .in0(N__38121),
            .in1(N__38112),
            .in2(_gnd_net_),
            .in3(N__38431),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_15_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_15_16_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_15_16_3  (
            .in0(N__47623),
            .in1(N__48243),
            .in2(N__42248),
            .in3(N__43256),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_15_16_5 .LUT_INIT=16'b0010011100100111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_15_16_5  (
            .in0(N__38432),
            .in1(N__38076),
            .in2(N__38067),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_16_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_16_6  (
            .in0(N__38040),
            .in1(N__38031),
            .in2(_gnd_net_),
            .in3(N__38429),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_15_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_15_16_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_15_16_7  (
            .in0(N__47619),
            .in1(N__48244),
            .in2(N__43163),
            .in3(N__42176),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_17_0 .LUT_INIT=16'b1111001111110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_17_0  (
            .in0(N__38276),
            .in1(N__48228),
            .in2(N__42318),
            .in3(N__47863),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_2  (
            .in0(N__48235),
            .in1(N__47862),
            .in2(N__42960),
            .in3(N__42458),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_3  (
            .in0(N__48227),
            .in1(N__40220),
            .in2(N__47879),
            .in3(N__42515),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_17_4 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_17_4  (
            .in0(N__43484),
            .in1(N__48225),
            .in2(N__43452),
            .in3(N__47857),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_17_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_17_5  (
            .in0(N__48226),
            .in1(N__42085),
            .in2(N__47878),
            .in3(N__40325),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_7  (
            .in0(N__47861),
            .in1(N__48234),
            .in2(N__43209),
            .in3(N__42657),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_18_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_18_1  (
            .in0(N__47848),
            .in1(N__48236),
            .in2(N__42912),
            .in3(N__42418),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_18_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_18_2  (
            .in0(N__48237),
            .in1(N__47849),
            .in2(N__43533),
            .in3(N__42352),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40008),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_15_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_15_19_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_15_19_5  (
            .in0(N__41575),
            .in1(N__41559),
            .in2(_gnd_net_),
            .in3(N__46955),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_15_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_15_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40203),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__38249),
            .in2(N__46554),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__38803),
            .in2(N__48486),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__39477),
            .in2(N__38849),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__38807),
            .in2(N__39816),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__39762),
            .in2(N__38850),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__38811),
            .in2(N__39711),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__39801),
            .in2(N__38851),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__38815),
            .in2(N__39492),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__38693),
            .in2(N__39888),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__39828),
            .in2(N__38749),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__38681),
            .in2(N__39843),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__43314),
            .in2(N__38746),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__38685),
            .in2(N__39981),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__43392),
            .in2(N__38747),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_22_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__38689),
            .in2(N__43407),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_22_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(N__39726),
            .in2(N__38748),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__39870),
            .in2(N__38759),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_23_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__38724),
            .in2(N__40518),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_23_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__40332),
            .in2(N__38760),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_23_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__38728),
            .in2(N__40347),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_23_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__40107),
            .in2(N__38761),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_23_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__38732),
            .in2(N__40293),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_23_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__39858),
            .in2(N__38762),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__38736),
            .in2(N__39924),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__38816),
            .in2(N__39954),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__40500),
            .in2(N__38852),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__38820),
            .in2(N__40284),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__40338),
            .in2(N__38853),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_24_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__38824),
            .in2(N__40494),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_24_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__40485),
            .in2(N__38854),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_24_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_15_24_6  (
            .in0(_gnd_net_),
            .in1(N__38828),
            .in2(N__40509),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_24_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_24_7  (
            .in0(N__48242),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38502),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_16_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_16_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_16_5_3 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_16_5_3  (
            .in0(N__38316),
            .in1(N__39060),
            .in2(N__39027),
            .in3(N__39372),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49942),
            .ce(),
            .sr(N__49293));
    defparam \phase_controller_inst2.stoper_hc.running_LC_16_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_16_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_16_5_5 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_16_5_5  (
            .in0(N__38292),
            .in1(N__39059),
            .in2(N__39026),
            .in3(N__39371),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49942),
            .ce(),
            .sr(N__49293));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_16_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_16_6_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__39018),
            .in2(_gnd_net_),
            .in3(N__39370),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38280),
            .in3(N__39061),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_6_2 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_6_2  (
            .in0(N__39063),
            .in1(N__41215),
            .in2(N__39039),
            .in3(N__40418),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(),
            .sr(N__49298));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_16_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_16_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_16_6_3  (
            .in0(_gnd_net_),
            .in1(N__39062),
            .in2(_gnd_net_),
            .in3(N__39035),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_6_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_6_7  (
            .in0(N__39019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38985),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_16_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_16_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(N__45117),
            .in2(N__38949),
            .in3(N__40414),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_16_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_16_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_16_7_1  (
            .in0(N__40397),
            .in1(N__38937),
            .in2(N__38931),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_16_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_16_7_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_16_7_2  (
            .in0(N__40373),
            .in1(N__38922),
            .in2(N__38916),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_16_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_16_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(N__38904),
            .in2(N__38898),
            .in3(N__40682),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_16_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_16_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__38889),
            .in2(N__38883),
            .in3(N__40667),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_16_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_16_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(N__45396),
            .in2(N__38871),
            .in3(N__40652),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_16_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_16_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(N__45321),
            .in2(N__39147),
            .in3(N__40637),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_16_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_16_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(N__39138),
            .in2(N__39123),
            .in3(N__40622),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_16_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_16_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_16_8_0  (
            .in0(N__40607),
            .in1(N__40881),
            .in2(N__39114),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_16_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_16_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__40971),
            .in2(N__39105),
            .in3(N__40592),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_16_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_16_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__39096),
            .in2(N__40905),
            .in3(N__40577),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_16_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_16_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__40893),
            .in2(N__39090),
            .in3(N__40802),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_16_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_16_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__45225),
            .in2(N__39081),
            .in3(N__40787),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_16_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_16_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_16_8_5  (
            .in0(N__40772),
            .in1(N__44502),
            .in2(N__39072),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_16_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_16_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__39228),
            .in2(N__45159),
            .in3(N__40757),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_16_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_16_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__44490),
            .in2(N__44433),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_16_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_16_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__39222),
            .in2(N__39210),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_16_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_16_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__44889),
            .in2(N__45531),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_16_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_16_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__41037),
            .in2(N__41097),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_16_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_16_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__45105),
            .in2(N__45051),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_16_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_16_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__44898),
            .in2(N__44961),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_16_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_16_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__39201),
            .in2(N__39186),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_16_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_16_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__39171),
            .in2(N__39162),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39375),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__45272),
            .in2(N__50355),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49885),
            .ce(N__50238),
            .sr(N__49329));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__45248),
            .in2(N__45306),
            .in3(N__39321),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49885),
            .ce(N__50238),
            .sr(N__49329));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__45273),
            .in2(N__45815),
            .in3(N__39282),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49885),
            .ce(N__50238),
            .sr(N__49329));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__45249),
            .in2(N__45785),
            .in3(N__39279),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49885),
            .ce(N__50238),
            .sr(N__49329));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__45755),
            .in2(N__45816),
            .in3(N__39276),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49885),
            .ce(N__50238),
            .sr(N__49329));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__45731),
            .in2(N__45786),
            .in3(N__39234),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49885),
            .ce(N__50238),
            .sr(N__49329));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__45756),
            .in2(N__45707),
            .in3(N__39231),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49885),
            .ce(N__50238),
            .sr(N__49329));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__45732),
            .in2(N__45668),
            .in3(N__39402),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49885),
            .ce(N__50238),
            .sr(N__49329));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__45626),
            .in2(N__45708),
            .in3(N__39399),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49875),
            .ce(N__50233),
            .sr(N__49337));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__45599),
            .in2(N__45669),
            .in3(N__39396),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49875),
            .ce(N__50233),
            .sr(N__49337));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__46085),
            .in2(N__45630),
            .in3(N__39393),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49875),
            .ce(N__50233),
            .sr(N__49337));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__45600),
            .in2(N__46058),
            .in3(N__39390),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49875),
            .ce(N__50233),
            .sr(N__49337));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__46025),
            .in2(N__46089),
            .in3(N__39387),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49875),
            .ce(N__50233),
            .sr(N__49337));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__45998),
            .in2(N__46059),
            .in3(N__39384),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49875),
            .ce(N__50233),
            .sr(N__49337));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__45971),
            .in2(N__46029),
            .in3(N__39381),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49875),
            .ce(N__50233),
            .sr(N__49337));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__45999),
            .in2(N__45938),
            .in3(N__39378),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49875),
            .ce(N__50233),
            .sr(N__49337));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__45902),
            .in2(N__45975),
            .in3(N__39429),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49864),
            .ce(N__50234),
            .sr(N__49346));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__45872),
            .in2(N__45939),
            .in3(N__39426),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49864),
            .ce(N__50234),
            .sr(N__49346));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__45842),
            .in2(N__45906),
            .in3(N__39423),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49864),
            .ce(N__50234),
            .sr(N__49346));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__46322),
            .in2(N__45876),
            .in3(N__39420),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49864),
            .ce(N__50234),
            .sr(N__49346));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(N__46292),
            .in2(N__45846),
            .in3(N__39417),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49864),
            .ce(N__50234),
            .sr(N__49346));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__46265),
            .in2(N__46326),
            .in3(N__39414),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49864),
            .ce(N__50234),
            .sr(N__49346));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(N__46238),
            .in2(N__46296),
            .in3(N__39411),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49864),
            .ce(N__50234),
            .sr(N__49346));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(N__46266),
            .in2(N__46205),
            .in3(N__39408),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49864),
            .ce(N__50234),
            .sr(N__49346));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__46166),
            .in2(N__46242),
            .in3(N__39405),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49853),
            .ce(N__50226),
            .sr(N__49356));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__46139),
            .in2(N__46206),
            .in3(N__39657),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49853),
            .ce(N__50226),
            .sr(N__49356));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__46167),
            .in2(N__46113),
            .in3(N__39615),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49853),
            .ce(N__50226),
            .sr(N__49356));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__46608),
            .in2(N__46143),
            .in3(N__39573),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49853),
            .ce(N__50226),
            .sr(N__49356));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39570),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(N__50226),
            .sr(N__49356));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_13_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__45305),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(N__50226),
            .sr(N__49356));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_16_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_16_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_16_14_1  (
            .in0(N__48087),
            .in1(N__42859),
            .in2(N__47875),
            .in3(N__41744),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46529),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49841),
            .ce(N__46411),
            .sr(N__49363));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_0  (
            .in0(N__40027),
            .in1(N__48584),
            .in2(_gnd_net_),
            .in3(N__41995),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_1  (
            .in0(N__48580),
            .in1(N__40081),
            .in2(_gnd_net_),
            .in3(N__41767),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_2  (
            .in0(N__42866),
            .in1(N__48581),
            .in2(_gnd_net_),
            .in3(N__41743),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_3  (
            .in0(N__48583),
            .in1(_gnd_net_),
            .in2(N__42757),
            .in3(N__42040),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_15_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_15_4  (
            .in0(N__47801),
            .in1(N__48091),
            .in2(N__42278),
            .in3(N__43103),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_15_5 .LUT_INIT=16'b1010001110100011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_15_5  (
            .in0(N__41717),
            .in1(N__41837),
            .in2(N__48198),
            .in3(N__47799),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_6  (
            .in0(N__41836),
            .in1(N__48582),
            .in2(_gnd_net_),
            .in3(N__41716),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_16_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_16_15_7 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_16_15_7  (
            .in0(N__42819),
            .in1(N__47800),
            .in2(N__41700),
            .in3(N__48092),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_16_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_16_0  (
            .in0(N__48186),
            .in1(N__47796),
            .in2(N__40166),
            .in3(N__41936),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_1  (
            .in0(N__43102),
            .in1(N__48624),
            .in2(_gnd_net_),
            .in3(N__42268),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_2  (
            .in0(N__48622),
            .in1(_gnd_net_),
            .in2(N__42817),
            .in3(N__41695),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_16_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_16_16_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_16_16_3  (
            .in0(N__47798),
            .in1(N__48187),
            .in2(N__47918),
            .in3(N__47272),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40080),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41827),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_16_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_16_6  (
            .in0(N__48185),
            .in1(N__47797),
            .in2(N__42818),
            .in3(N__41696),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_7  (
            .in0(N__42697),
            .in1(N__48623),
            .in2(_gnd_net_),
            .in3(N__41965),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_0  (
            .in0(N__48628),
            .in1(N__43249),
            .in2(_gnd_net_),
            .in3(N__42235),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_1  (
            .in0(N__48638),
            .in1(N__40256),
            .in2(_gnd_net_),
            .in3(N__42550),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_17_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_17_2  (
            .in0(N__48626),
            .in1(N__48352),
            .in2(_gnd_net_),
            .in3(N__48385),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_17_3 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_17_3  (
            .in0(N__40159),
            .in1(N__41935),
            .in2(_gnd_net_),
            .in3(N__48625),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40158),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_17_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_17_5  (
            .in0(N__48460),
            .in1(N__48627),
            .in2(_gnd_net_),
            .in3(N__48421),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48384),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43371),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40317),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_1  (
            .in0(N__40249),
            .in1(N__48197),
            .in2(N__47877),
            .in3(N__42551),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40548),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_3  (
            .in0(N__48640),
            .in1(N__43048),
            .in2(_gnd_net_),
            .in3(N__42478),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_18_4 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_18_4  (
            .in0(N__48196),
            .in1(N__47853),
            .in2(N__48291),
            .in3(N__48314),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_5  (
            .in0(N__48639),
            .in1(N__40213),
            .in2(_gnd_net_),
            .in3(N__42508),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_6  (
            .in0(N__48644),
            .in1(N__48313),
            .in2(_gnd_net_),
            .in3(N__48286),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_18_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_18_7  (
            .in0(N__40248),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__46490),
            .in2(N__43299),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49816),
            .ce(N__46410),
            .sr(N__49388));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__46439),
            .in2(N__43805),
            .in3(N__40053),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49816),
            .ce(N__46410),
            .sr(N__49388));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__43298),
            .in2(N__43775),
            .in3(N__40050),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49816),
            .ce(N__46410),
            .sr(N__49388));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__43742),
            .in2(N__43806),
            .in3(N__40047),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49816),
            .ce(N__46410),
            .sr(N__49388));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__43715),
            .in2(N__43776),
            .in3(N__40044),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49816),
            .ce(N__46410),
            .sr(N__49388));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__43691),
            .in2(N__43746),
            .in3(N__39987),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49816),
            .ce(N__46410),
            .sr(N__49388));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__43716),
            .in2(N__43667),
            .in3(N__39984),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49816),
            .ce(N__46410),
            .sr(N__49388));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__43692),
            .in2(N__43635),
            .in3(N__40134),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49816),
            .ce(N__46410),
            .sr(N__49388));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__43592),
            .in2(N__43668),
            .in3(N__40131),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49815),
            .ce(N__46409),
            .sr(N__49392));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__43565),
            .in2(N__43634),
            .in3(N__40128),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49815),
            .ce(N__46409),
            .sr(N__49392));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__44033),
            .in2(N__43596),
            .in3(N__40125),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49815),
            .ce(N__46409),
            .sr(N__49392));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__43566),
            .in2(N__44009),
            .in3(N__40122),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49815),
            .ce(N__46409),
            .sr(N__49392));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__44034),
            .in2(N__43979),
            .in3(N__40119),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49815),
            .ce(N__46409),
            .sr(N__49392));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(N__43946),
            .in2(N__44010),
            .in3(N__40116),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49815),
            .ce(N__46409),
            .sr(N__49392));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__43916),
            .in2(N__43980),
            .in3(N__40113),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49815),
            .ce(N__46409),
            .sr(N__49392));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__43886),
            .in2(N__43950),
            .in3(N__40110),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49815),
            .ce(N__46409),
            .sr(N__49392));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__43853),
            .in2(N__43920),
            .in3(N__40275),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49813),
            .ce(N__46408),
            .sr(N__49396));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__43829),
            .in2(N__43890),
            .in3(N__40272),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49813),
            .ce(N__46408),
            .sr(N__49396));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__43854),
            .in2(N__44288),
            .in3(N__40269),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49813),
            .ce(N__46408),
            .sr(N__49396));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__43830),
            .in2(N__44258),
            .in3(N__40266),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49813),
            .ce(N__46408),
            .sr(N__49396));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__44228),
            .in2(N__44289),
            .in3(N__40224),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49813),
            .ce(N__46408),
            .sr(N__49396));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(N__44201),
            .in2(N__44259),
            .in3(N__40182),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49813),
            .ce(N__46408),
            .sr(N__49396));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(N__44229),
            .in2(N__44174),
            .in3(N__40179),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49813),
            .ce(N__46408),
            .sr(N__49396));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(N__44138),
            .in2(N__44205),
            .in3(N__40176),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49813),
            .ce(N__46408),
            .sr(N__49396));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__44102),
            .in2(N__44175),
            .in3(N__40173),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49811),
            .ce(N__46407),
            .sr(N__49399));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(N__44075),
            .in2(N__44142),
            .in3(N__40359),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49811),
            .ce(N__46407),
            .sr(N__49399));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(N__44052),
            .in2(N__44106),
            .in3(N__40356),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49811),
            .ce(N__46407),
            .sr(N__49399));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__44076),
            .in2(N__44736),
            .in3(N__40353),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49811),
            .ce(N__46407),
            .sr(N__49399));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40350),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_23_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_23_0  (
            .in0(N__42598),
            .in1(N__48647),
            .in2(_gnd_net_),
            .in3(N__42136),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_1  (
            .in0(N__42896),
            .in1(N__48184),
            .in2(_gnd_net_),
            .in3(N__42420),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_23_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_23_3  (
            .in0(N__48646),
            .in1(N__43150),
            .in2(_gnd_net_),
            .in3(N__42175),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_23_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_23_4  (
            .in0(N__40324),
            .in1(N__48648),
            .in2(_gnd_net_),
            .in3(N__42089),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_5  (
            .in0(N__42940),
            .in1(N__48183),
            .in2(_gnd_net_),
            .in3(N__42459),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_23_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_23_7  (
            .in0(N__48645),
            .in1(N__40552),
            .in2(_gnd_net_),
            .in3(N__42212),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_24_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(N__48182),
            .in2(_gnd_net_),
            .in3(N__42314),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_24_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_24_2  (
            .in0(N__48179),
            .in1(N__43201),
            .in2(_gnd_net_),
            .in3(N__42656),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_24_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_24_4  (
            .in0(N__48180),
            .in1(N__42997),
            .in2(_gnd_net_),
            .in3(N__42388),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_24_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_24_7  (
            .in0(N__43519),
            .in1(N__48181),
            .in2(_gnd_net_),
            .in3(N__42354),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_17_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_17_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_17_6_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_17_6_2  (
            .in0(N__40479),
            .in1(N__47047),
            .in2(_gnd_net_),
            .in3(N__40440),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(N__47160),
            .sr(N__49294));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(N__40425),
            .in2(N__40419),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_7_1  (
            .in0(N__41211),
            .in1(N__40398),
            .in2(_gnd_net_),
            .in3(N__40386),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49933),
            .ce(),
            .sr(N__49299));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_7_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_7_2  (
            .in0(N__41263),
            .in1(N__40374),
            .in2(N__40383),
            .in3(N__40362),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49933),
            .ce(),
            .sr(N__49299));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_7_3  (
            .in0(N__41212),
            .in1(N__40683),
            .in2(_gnd_net_),
            .in3(N__40671),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49933),
            .ce(),
            .sr(N__49299));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_7_4  (
            .in0(N__41264),
            .in1(N__40668),
            .in2(_gnd_net_),
            .in3(N__40656),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49933),
            .ce(),
            .sr(N__49299));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_7_5  (
            .in0(N__41213),
            .in1(N__40653),
            .in2(_gnd_net_),
            .in3(N__40641),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49933),
            .ce(),
            .sr(N__49299));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_7_6  (
            .in0(N__41265),
            .in1(N__40638),
            .in2(_gnd_net_),
            .in3(N__40626),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49933),
            .ce(),
            .sr(N__49299));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_7_7  (
            .in0(N__41214),
            .in1(N__40623),
            .in2(_gnd_net_),
            .in3(N__40611),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49933),
            .ce(),
            .sr(N__49299));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_8_0  (
            .in0(N__41253),
            .in1(N__40608),
            .in2(_gnd_net_),
            .in3(N__40596),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49921),
            .ce(),
            .sr(N__49307));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_8_1  (
            .in0(N__41242),
            .in1(N__40593),
            .in2(_gnd_net_),
            .in3(N__40581),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49921),
            .ce(),
            .sr(N__49307));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_8_2  (
            .in0(N__41250),
            .in1(N__40578),
            .in2(_gnd_net_),
            .in3(N__40566),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49921),
            .ce(),
            .sr(N__49307));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_8_3  (
            .in0(N__41243),
            .in1(N__40803),
            .in2(_gnd_net_),
            .in3(N__40791),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49921),
            .ce(),
            .sr(N__49307));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_8_4  (
            .in0(N__41251),
            .in1(N__40788),
            .in2(_gnd_net_),
            .in3(N__40776),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49921),
            .ce(),
            .sr(N__49307));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_8_5  (
            .in0(N__41244),
            .in1(N__40773),
            .in2(_gnd_net_),
            .in3(N__40761),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49921),
            .ce(),
            .sr(N__49307));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_8_6  (
            .in0(N__41252),
            .in1(N__40758),
            .in2(_gnd_net_),
            .in3(N__40746),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49921),
            .ce(),
            .sr(N__49307));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_8_7  (
            .in0(N__41245),
            .in1(N__44477),
            .in2(_gnd_net_),
            .in3(N__40743),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49921),
            .ce(),
            .sr(N__49307));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_9_0  (
            .in0(N__41246),
            .in1(N__44459),
            .in2(_gnd_net_),
            .in3(N__40740),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_9_1  (
            .in0(N__41276),
            .in1(N__40727),
            .in2(_gnd_net_),
            .in3(N__40713),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_9_2  (
            .in0(N__41247),
            .in1(N__40703),
            .in2(_gnd_net_),
            .in3(N__40689),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_9_3  (
            .in0(N__41277),
            .in1(N__45546),
            .in2(_gnd_net_),
            .in3(N__40686),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_9_4  (
            .in0(N__41248),
            .in1(N__45563),
            .in2(_gnd_net_),
            .in3(N__40869),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_9_5  (
            .in0(N__41278),
            .in1(N__41056),
            .in2(_gnd_net_),
            .in3(N__40866),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_9_6  (
            .in0(N__41249),
            .in1(N__41077),
            .in2(_gnd_net_),
            .in3(N__40863),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_9_7  (
            .in0(N__41279),
            .in1(N__45066),
            .in2(_gnd_net_),
            .in3(N__40860),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49910),
            .ce(),
            .sr(N__49314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_10_0  (
            .in0(N__41269),
            .in1(N__45083),
            .in2(_gnd_net_),
            .in3(N__40857),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49899),
            .ce(),
            .sr(N__49321));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_10_1  (
            .in0(N__41273),
            .in1(N__44948),
            .in2(_gnd_net_),
            .in3(N__40854),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49899),
            .ce(),
            .sr(N__49321));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_10_2  (
            .in0(N__41270),
            .in1(N__44916),
            .in2(_gnd_net_),
            .in3(N__40851),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49899),
            .ce(),
            .sr(N__49321));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_10_3  (
            .in0(N__41274),
            .in1(N__40846),
            .in2(_gnd_net_),
            .in3(N__40830),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49899),
            .ce(),
            .sr(N__49321));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_10_4  (
            .in0(N__41271),
            .in1(N__40822),
            .in2(_gnd_net_),
            .in3(N__40806),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49899),
            .ce(),
            .sr(N__49321));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_10_5  (
            .in0(N__41275),
            .in1(N__41308),
            .in2(_gnd_net_),
            .in3(N__41289),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49899),
            .ce(),
            .sr(N__49321));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_10_6  (
            .in0(N__41272),
            .in1(N__41119),
            .in2(_gnd_net_),
            .in3(N__41130),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49899),
            .ce(),
            .sr(N__49321));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_11_0 .LUT_INIT=16'b0100111100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_11_0  (
            .in0(N__41057),
            .in1(N__41640),
            .in2(N__41082),
            .in3(N__41526),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_17_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_17_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_17_11_1  (
            .in0(N__41639),
            .in1(N__41081),
            .in2(N__41061),
            .in3(N__41525),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_17_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_17_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_17_11_4  (
            .in0(N__41028),
            .in1(N__40987),
            .in2(_gnd_net_),
            .in3(N__47021),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49886),
            .ce(N__47155),
            .sr(N__49330));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_17_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_17_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_17_11_5  (
            .in0(N__47020),
            .in1(N__40947),
            .in2(_gnd_net_),
            .in3(N__40929),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49886),
            .ce(N__47155),
            .sr(N__49330));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_17_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_17_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_17_11_6  (
            .in0(N__41367),
            .in1(N__41342),
            .in2(_gnd_net_),
            .in3(N__47022),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49886),
            .ce(N__47155),
            .sr(N__49330));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_17_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_17_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_17_12_0  (
            .in0(N__47024),
            .in1(N__41395),
            .in2(_gnd_net_),
            .in3(N__41431),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(N__47154),
            .sr(N__49338));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_17_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_17_12_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_17_12_1  (
            .in0(N__41678),
            .in1(N__47025),
            .in2(_gnd_net_),
            .in3(N__41655),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(N__47154),
            .sr(N__49338));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_17_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_17_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_17_12_4  (
            .in0(N__47023),
            .in1(N__41623),
            .in2(_gnd_net_),
            .in3(N__41604),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(N__47154),
            .sr(N__49338));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_17_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_17_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_17_12_5  (
            .in0(N__41586),
            .in1(N__41551),
            .in2(_gnd_net_),
            .in3(N__47026),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49876),
            .ce(N__47154),
            .sr(N__49338));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_17_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_17_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_17_13_0  (
            .in0(N__46874),
            .in1(N__41461),
            .in2(_gnd_net_),
            .in3(N__41513),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_13_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_13_2  (
            .in0(N__46464),
            .in1(N__48086),
            .in2(_gnd_net_),
            .in3(N__41892),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_13_3  (
            .in0(N__44347),
            .in1(N__44320),
            .in2(_gnd_net_),
            .in3(N__46875),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_17_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_17_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_17_13_5  (
            .in0(N__45139),
            .in1(N__46880),
            .in2(_gnd_net_),
            .in3(N__50324),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_13_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_13_6  (
            .in0(N__41430),
            .in1(_gnd_net_),
            .in2(N__46991),
            .in3(N__41396),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_13_7  (
            .in0(N__41341),
            .in1(N__41374),
            .in2(_gnd_net_),
            .in3(N__46879),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46577),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_14_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__48008),
            .in2(N__41886),
            .in3(N__46460),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_17_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_17_14_3 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_17_14_3  (
            .in0(N__48507),
            .in1(N__48524),
            .in2(N__46376),
            .in3(N__48009),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_6  (
            .in0(N__48010),
            .in1(N__41838),
            .in2(N__47876),
            .in3(N__41718),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__46383),
            .in2(N__46578),
            .in3(N__46576),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__41787),
            .in2(_gnd_net_),
            .in3(N__41754),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__42828),
            .in2(_gnd_net_),
            .in3(N__41727),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__41724),
            .in2(_gnd_net_),
            .in3(N__41703),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__42786),
            .in2(_gnd_net_),
            .in3(N__42057),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__42723),
            .in2(_gnd_net_),
            .in3(N__42024),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__42021),
            .in2(_gnd_net_),
            .in3(N__41979),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__42669),
            .in2(_gnd_net_),
            .in3(N__41952),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__41949),
            .in2(_gnd_net_),
            .in3(N__41919),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__41916),
            .in2(_gnd_net_),
            .in3(N__41910),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__41907),
            .in2(_gnd_net_),
            .in3(N__41901),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__42768),
            .in2(_gnd_net_),
            .in3(N__41898),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__42777),
            .in2(_gnd_net_),
            .in3(N__41895),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__43269),
            .in2(_gnd_net_),
            .in3(N__42282),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__43074),
            .in2(_gnd_net_),
            .in3(N__42252),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__43218),
            .in2(_gnd_net_),
            .in3(N__42222),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__42219),
            .in2(_gnd_net_),
            .in3(N__42183),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43122),
            .in3(N__42144),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__42573),
            .in2(_gnd_net_),
            .in3(N__42105),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__43542),
            .in2(_gnd_net_),
            .in3(N__42102),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__42099),
            .in2(_gnd_net_),
            .in3(N__42060),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__42564),
            .in2(_gnd_net_),
            .in3(N__42534),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__42531),
            .in2(_gnd_net_),
            .in3(N__42492),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__43023),
            .in2(_gnd_net_),
            .in3(N__42465),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__43173),
            .in2(_gnd_net_),
            .in3(N__42462),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__42921),
            .in2(_gnd_net_),
            .in3(N__42423),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__42879),
            .in2(_gnd_net_),
            .in3(N__42393),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__42969),
            .in2(_gnd_net_),
            .in3(N__42357),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__43494),
            .in2(_gnd_net_),
            .in3(N__42324),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42321),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_18_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_18_6  (
            .in0(N__42844),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42799),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47901),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48450),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42738),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42687),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_19_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_19_7  (
            .in0(N__48254),
            .in1(N__42640),
            .in2(N__47880),
            .in3(N__43205),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42589),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43470),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43239),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43191),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43140),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43092),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43039),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42987),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42939),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42895),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48304),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43510),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_22_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_22_1  (
            .in0(N__48643),
            .in1(N__43480),
            .in2(_gnd_net_),
            .in3(N__43441),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_22_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_22_2  (
            .in0(N__47911),
            .in1(N__48642),
            .in2(_gnd_net_),
            .in3(N__47277),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_22_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_22_3  (
            .in0(N__48641),
            .in1(N__43375),
            .in2(_gnd_net_),
            .in3(N__43336),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_17_23_0  (
            .in0(N__44867),
            .in1(N__46483),
            .in2(_gnd_net_),
            .in3(N__43305),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__49812),
            .ce(N__44714),
            .sr(N__49400));
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_17_23_1  (
            .in0(N__44818),
            .in1(N__46432),
            .in2(_gnd_net_),
            .in3(N__43302),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__49812),
            .ce(N__44714),
            .sr(N__49400));
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_17_23_2  (
            .in0(N__44868),
            .in1(N__43288),
            .in2(_gnd_net_),
            .in3(N__43272),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__49812),
            .ce(N__44714),
            .sr(N__49400));
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_17_23_3  (
            .in0(N__44819),
            .in1(N__43793),
            .in2(_gnd_net_),
            .in3(N__43779),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__49812),
            .ce(N__44714),
            .sr(N__49400));
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_17_23_4  (
            .in0(N__44869),
            .in1(N__43763),
            .in2(_gnd_net_),
            .in3(N__43749),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__49812),
            .ce(N__44714),
            .sr(N__49400));
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_17_23_5  (
            .in0(N__44820),
            .in1(N__43735),
            .in2(_gnd_net_),
            .in3(N__43719),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__49812),
            .ce(N__44714),
            .sr(N__49400));
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_17_23_6  (
            .in0(N__44870),
            .in1(N__43709),
            .in2(_gnd_net_),
            .in3(N__43695),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__49812),
            .ce(N__44714),
            .sr(N__49400));
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_17_23_7  (
            .in0(N__44821),
            .in1(N__43685),
            .in2(_gnd_net_),
            .in3(N__43671),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__49812),
            .ce(N__44714),
            .sr(N__49400));
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_17_24_0  (
            .in0(N__44849),
            .in1(N__43654),
            .in2(_gnd_net_),
            .in3(N__43638),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__49810),
            .ce(N__44706),
            .sr(N__49406));
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_17_24_1  (
            .in0(N__44853),
            .in1(N__43618),
            .in2(_gnd_net_),
            .in3(N__43599),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__49810),
            .ce(N__44706),
            .sr(N__49406));
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_17_24_2  (
            .in0(N__44846),
            .in1(N__43585),
            .in2(_gnd_net_),
            .in3(N__43569),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__49810),
            .ce(N__44706),
            .sr(N__49406));
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_17_24_3  (
            .in0(N__44850),
            .in1(N__43559),
            .in2(_gnd_net_),
            .in3(N__43545),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__49810),
            .ce(N__44706),
            .sr(N__49406));
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_17_24_4  (
            .in0(N__44847),
            .in1(N__44027),
            .in2(_gnd_net_),
            .in3(N__44013),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__49810),
            .ce(N__44706),
            .sr(N__49406));
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_17_24_5  (
            .in0(N__44851),
            .in1(N__43997),
            .in2(_gnd_net_),
            .in3(N__43983),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__49810),
            .ce(N__44706),
            .sr(N__49406));
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_17_24_6  (
            .in0(N__44848),
            .in1(N__43967),
            .in2(_gnd_net_),
            .in3(N__43953),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__49810),
            .ce(N__44706),
            .sr(N__49406));
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_17_24_7  (
            .in0(N__44852),
            .in1(N__43939),
            .in2(_gnd_net_),
            .in3(N__43923),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__49810),
            .ce(N__44706),
            .sr(N__49406));
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_17_25_0  (
            .in0(N__44863),
            .in1(N__43909),
            .in2(_gnd_net_),
            .in3(N__43893),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_25_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__49807),
            .ce(N__44715),
            .sr(N__49409));
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_17_25_1  (
            .in0(N__44871),
            .in1(N__43879),
            .in2(_gnd_net_),
            .in3(N__43857),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__49807),
            .ce(N__44715),
            .sr(N__49409));
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_17_25_2  (
            .in0(N__44864),
            .in1(N__43847),
            .in2(_gnd_net_),
            .in3(N__43833),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__49807),
            .ce(N__44715),
            .sr(N__49409));
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_17_25_3  (
            .in0(N__44872),
            .in1(N__43823),
            .in2(_gnd_net_),
            .in3(N__43809),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__49807),
            .ce(N__44715),
            .sr(N__49409));
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_17_25_4  (
            .in0(N__44865),
            .in1(N__44276),
            .in2(_gnd_net_),
            .in3(N__44262),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__49807),
            .ce(N__44715),
            .sr(N__49409));
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_25_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_17_25_5  (
            .in0(N__44873),
            .in1(N__44246),
            .in2(_gnd_net_),
            .in3(N__44232),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__49807),
            .ce(N__44715),
            .sr(N__49409));
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_25_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_17_25_6  (
            .in0(N__44866),
            .in1(N__44222),
            .in2(_gnd_net_),
            .in3(N__44208),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__49807),
            .ce(N__44715),
            .sr(N__49409));
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_25_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_17_25_7  (
            .in0(N__44874),
            .in1(N__44194),
            .in2(_gnd_net_),
            .in3(N__44178),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__49807),
            .ce(N__44715),
            .sr(N__49409));
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_26_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_17_26_0  (
            .in0(N__44822),
            .in1(N__44161),
            .in2(_gnd_net_),
            .in3(N__44145),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_26_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__49804),
            .ce(N__44713),
            .sr(N__49413));
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_26_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_26_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_17_26_1  (
            .in0(N__44826),
            .in1(N__44131),
            .in2(_gnd_net_),
            .in3(N__44109),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__49804),
            .ce(N__44713),
            .sr(N__49413));
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_26_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_17_26_2  (
            .in0(N__44823),
            .in1(N__44095),
            .in2(_gnd_net_),
            .in3(N__44079),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__49804),
            .ce(N__44713),
            .sr(N__49413));
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_26_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_17_26_3  (
            .in0(N__44827),
            .in1(N__44069),
            .in2(_gnd_net_),
            .in3(N__44055),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__49804),
            .ce(N__44713),
            .sr(N__49413));
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_26_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_26_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_17_26_4  (
            .in0(N__44824),
            .in1(N__44048),
            .in2(_gnd_net_),
            .in3(N__44877),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__49804),
            .ce(N__44713),
            .sr(N__49413));
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_26_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_26_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_17_26_5  (
            .in0(N__44729),
            .in1(N__44825),
            .in2(_gnd_net_),
            .in3(N__44739),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(N__44713),
            .sr(N__49413));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_18_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_18_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_18_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_18_7_0  (
            .in0(N__47040),
            .in1(N__44667),
            .in2(_gnd_net_),
            .in3(N__44631),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49944),
            .ce(N__47161),
            .sr(N__49295));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_18_7_5  (
            .in0(N__44613),
            .in1(N__44588),
            .in2(_gnd_net_),
            .in3(N__47042),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49944),
            .ce(N__47161),
            .sr(N__49295));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_18_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_18_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_18_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_18_7_7  (
            .in0(N__44547),
            .in1(N__44517),
            .in2(_gnd_net_),
            .in3(N__47041),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49944),
            .ce(N__47161),
            .sr(N__49295));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_8_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_8_0  (
            .in0(N__44442),
            .in1(N__44364),
            .in2(N__44478),
            .in3(N__44458),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_8_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_8_1  (
            .in0(N__44363),
            .in1(N__44476),
            .in2(N__44460),
            .in3(N__44441),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_18_8_2  (
            .in0(N__44418),
            .in1(N__47044),
            .in2(_gnd_net_),
            .in3(N__44382),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(N__47159),
            .sr(N__49300));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_18_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_18_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_18_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_18_8_4  (
            .in0(N__44355),
            .in1(N__44325),
            .in2(_gnd_net_),
            .in3(N__47045),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(N__47159),
            .sr(N__49300));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_18_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_18_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_18_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_18_8_6  (
            .in0(N__45216),
            .in1(N__45192),
            .in2(_gnd_net_),
            .in3(N__47046),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(N__47159),
            .sr(N__49300));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_18_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_18_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_18_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_18_8_7  (
            .in0(N__47043),
            .in1(N__45147),
            .in2(_gnd_net_),
            .in3(N__50323),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49934),
            .ce(N__47159),
            .sr(N__49300));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_9_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_9_0  (
            .in0(N__45065),
            .in1(N__45096),
            .in2(N__44973),
            .in3(N__45082),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_9_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_9_1  (
            .in0(N__45095),
            .in1(N__44972),
            .in2(N__45084),
            .in3(N__45064),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_18_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_18_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_18_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_18_9_3  (
            .in0(N__45039),
            .in1(N__45013),
            .in2(_gnd_net_),
            .in3(N__47032),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__47158),
            .sr(N__49308));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_9_5 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_9_5  (
            .in0(N__44927),
            .in1(N__44914),
            .in2(N__44949),
            .in3(N__47174),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_9_6 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_9_6  (
            .in0(N__44947),
            .in1(N__44928),
            .in2(N__47178),
            .in3(N__44915),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_10_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_10_0  (
            .in0(N__45545),
            .in1(N__45576),
            .in2(N__45456),
            .in3(N__45562),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_10_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_10_1  (
            .in0(N__45575),
            .in1(N__45455),
            .in2(N__45564),
            .in3(N__45544),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_18_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_18_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_18_10_3  (
            .in0(N__45515),
            .in1(N__47056),
            .in2(_gnd_net_),
            .in3(N__45474),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49911),
            .ce(N__47157),
            .sr(N__49315));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_18_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_18_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_18_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_18_10_4  (
            .in0(N__47055),
            .in1(N__45441),
            .in2(_gnd_net_),
            .in3(N__45414),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49911),
            .ce(N__47157),
            .sr(N__49315));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_18_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_18_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_18_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_18_10_5  (
            .in0(N__45384),
            .in1(N__47057),
            .in2(_gnd_net_),
            .in3(N__45352),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49911),
            .ce(N__47157),
            .sr(N__49315));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_11_0  (
            .in0(N__50177),
            .in1(N__50344),
            .in2(_gnd_net_),
            .in3(N__45309),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__49900),
            .ce(N__50283),
            .sr(N__49322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_11_1  (
            .in0(N__50173),
            .in1(N__45295),
            .in2(_gnd_net_),
            .in3(N__45276),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__49900),
            .ce(N__50283),
            .sr(N__49322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_11_2  (
            .in0(N__50178),
            .in1(N__45266),
            .in2(_gnd_net_),
            .in3(N__45252),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__49900),
            .ce(N__50283),
            .sr(N__49322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_11_3  (
            .in0(N__50174),
            .in1(N__45242),
            .in2(_gnd_net_),
            .in3(N__45228),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__49900),
            .ce(N__50283),
            .sr(N__49322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_11_4  (
            .in0(N__50179),
            .in1(N__45803),
            .in2(_gnd_net_),
            .in3(N__45789),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__49900),
            .ce(N__50283),
            .sr(N__49322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_11_5  (
            .in0(N__50175),
            .in1(N__45773),
            .in2(_gnd_net_),
            .in3(N__45759),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__49900),
            .ce(N__50283),
            .sr(N__49322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_11_6  (
            .in0(N__50180),
            .in1(N__45749),
            .in2(_gnd_net_),
            .in3(N__45735),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__49900),
            .ce(N__50283),
            .sr(N__49322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_11_7  (
            .in0(N__50176),
            .in1(N__45725),
            .in2(_gnd_net_),
            .in3(N__45711),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__49900),
            .ce(N__50283),
            .sr(N__49322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_12_0  (
            .in0(N__50166),
            .in1(N__45694),
            .in2(_gnd_net_),
            .in3(N__45672),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__49887),
            .ce(N__50278),
            .sr(N__49331));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_12_1  (
            .in0(N__50162),
            .in1(N__45655),
            .in2(_gnd_net_),
            .in3(N__45633),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__49887),
            .ce(N__50278),
            .sr(N__49331));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_12_2  (
            .in0(N__50163),
            .in1(N__45619),
            .in2(_gnd_net_),
            .in3(N__45603),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__49887),
            .ce(N__50278),
            .sr(N__49331));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_12_3  (
            .in0(N__50159),
            .in1(N__45593),
            .in2(_gnd_net_),
            .in3(N__45579),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__49887),
            .ce(N__50278),
            .sr(N__49331));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_12_4  (
            .in0(N__50164),
            .in1(N__46078),
            .in2(_gnd_net_),
            .in3(N__46062),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__49887),
            .ce(N__50278),
            .sr(N__49331));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_12_5  (
            .in0(N__50160),
            .in1(N__46046),
            .in2(_gnd_net_),
            .in3(N__46032),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__49887),
            .ce(N__50278),
            .sr(N__49331));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_12_6  (
            .in0(N__50165),
            .in1(N__46018),
            .in2(_gnd_net_),
            .in3(N__46002),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__49887),
            .ce(N__50278),
            .sr(N__49331));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_12_7  (
            .in0(N__50161),
            .in1(N__45997),
            .in2(_gnd_net_),
            .in3(N__45978),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__49887),
            .ce(N__50278),
            .sr(N__49331));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_13_0  (
            .in0(N__50146),
            .in1(N__45964),
            .in2(_gnd_net_),
            .in3(N__45942),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__49877),
            .ce(N__50277),
            .sr(N__49339));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_13_1  (
            .in0(N__50181),
            .in1(N__45925),
            .in2(_gnd_net_),
            .in3(N__45909),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__49877),
            .ce(N__50277),
            .sr(N__49339));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_13_2  (
            .in0(N__50147),
            .in1(N__45895),
            .in2(_gnd_net_),
            .in3(N__45879),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__49877),
            .ce(N__50277),
            .sr(N__49339));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_13_3  (
            .in0(N__50182),
            .in1(N__45865),
            .in2(_gnd_net_),
            .in3(N__45849),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__49877),
            .ce(N__50277),
            .sr(N__49339));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_13_4  (
            .in0(N__50148),
            .in1(N__45835),
            .in2(_gnd_net_),
            .in3(N__45819),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__49877),
            .ce(N__50277),
            .sr(N__49339));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_13_5  (
            .in0(N__50183),
            .in1(N__46315),
            .in2(_gnd_net_),
            .in3(N__46299),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__49877),
            .ce(N__50277),
            .sr(N__49339));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_13_6  (
            .in0(N__50149),
            .in1(N__46285),
            .in2(_gnd_net_),
            .in3(N__46269),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__49877),
            .ce(N__50277),
            .sr(N__49339));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_13_7  (
            .in0(N__50184),
            .in1(N__46259),
            .in2(_gnd_net_),
            .in3(N__46245),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__49877),
            .ce(N__50277),
            .sr(N__49339));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_14_0  (
            .in0(N__50167),
            .in1(N__46237),
            .in2(_gnd_net_),
            .in3(N__46209),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__49865),
            .ce(N__50279),
            .sr(N__49347));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_14_1  (
            .in0(N__50171),
            .in1(N__46192),
            .in2(_gnd_net_),
            .in3(N__46170),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__49865),
            .ce(N__50279),
            .sr(N__49347));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_14_2  (
            .in0(N__50168),
            .in1(N__46160),
            .in2(_gnd_net_),
            .in3(N__46146),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__49865),
            .ce(N__50279),
            .sr(N__49347));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_14_3  (
            .in0(N__50172),
            .in1(N__46132),
            .in2(_gnd_net_),
            .in3(N__46116),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__49865),
            .ce(N__50279),
            .sr(N__49347));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_14_4  (
            .in0(N__50169),
            .in1(N__46106),
            .in2(_gnd_net_),
            .in3(N__46092),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__49865),
            .ce(N__50279),
            .sr(N__49347));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_14_5  (
            .in0(N__46604),
            .in1(N__50170),
            .in2(_gnd_net_),
            .in3(N__46611),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49865),
            .ce(N__50279),
            .sr(N__49347));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_15_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__48206),
            .in2(_gnd_net_),
            .in3(N__47768),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46458),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_15_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_15_5  (
            .in0(N__46459),
            .in1(_gnd_net_),
            .in2(N__46557),
            .in3(N__48550),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46530),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(N__46413),
            .sr(N__49357));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46494),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(N__46413),
            .sr(N__49357));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46440),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49842),
            .ce(N__46412),
            .sr(N__49364));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48501),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3  (
            .in0(N__48503),
            .in1(N__48205),
            .in2(N__46377),
            .in3(N__48525),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4  (
            .in0(N__48551),
            .in1(N__48523),
            .in2(_gnd_net_),
            .in3(N__48502),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_18_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_18_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_18_17_1  (
            .in0(N__48239),
            .in1(N__48468),
            .in2(N__47865),
            .in3(N__48425),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_17_3  (
            .in0(N__48238),
            .in1(N__48392),
            .in2(N__47864),
            .in3(N__48353),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_18_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_18_17_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_18_17_5  (
            .in0(N__48241),
            .in1(N__47791),
            .in2(N__48321),
            .in3(N__48287),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_17_7  (
            .in0(N__48240),
            .in1(N__47919),
            .in2(N__47866),
            .in3(N__47273),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_20_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_20_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_20_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_20_8_7  (
            .in0(N__47244),
            .in1(N__47069),
            .in2(_gnd_net_),
            .in3(N__47211),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49949),
            .ce(N__47163),
            .sr(N__49301));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_20_9_4  (
            .in0(N__47120),
            .in1(N__50371),
            .in2(_gnd_net_),
            .in3(N__47070),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(N__47162),
            .sr(N__49309));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_20_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_20_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_20_10_5  (
            .in0(N__50375),
            .in1(N__47113),
            .in2(_gnd_net_),
            .in3(N__47048),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_20_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_20_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_20_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_20_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50351),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49923),
            .ce(N__50214),
            .sr(N__49323));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_20_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_20_13_4 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_20_13_4  (
            .in0(N__49972),
            .in1(_gnd_net_),
            .in2(N__50042),
            .in3(N__50006),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_164_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_20_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_20_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_20_13_5  (
            .in0(_gnd_net_),
            .in1(N__49973),
            .in2(_gnd_net_),
            .in3(N__50035),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_163_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_20_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_20_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_20_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49971),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_20_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_20_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_20_14_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_20_14_4  (
            .in0(N__49974),
            .in1(N__50043),
            .in2(_gnd_net_),
            .in3(N__50010),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49889),
            .ce(),
            .sr(N__49348));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_0  (
            .in0(N__48954),
            .in1(N__48881),
            .in2(_gnd_net_),
            .in3(N__48868),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
