// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 3 2024 21:46:45

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    error_pin,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    input error_pin;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__54407;
    wire N__54406;
    wire N__54405;
    wire N__54396;
    wire N__54395;
    wire N__54394;
    wire N__54387;
    wire N__54386;
    wire N__54385;
    wire N__54378;
    wire N__54377;
    wire N__54376;
    wire N__54369;
    wire N__54368;
    wire N__54367;
    wire N__54360;
    wire N__54359;
    wire N__54358;
    wire N__54351;
    wire N__54350;
    wire N__54349;
    wire N__54342;
    wire N__54341;
    wire N__54340;
    wire N__54333;
    wire N__54332;
    wire N__54331;
    wire N__54324;
    wire N__54323;
    wire N__54322;
    wire N__54315;
    wire N__54314;
    wire N__54313;
    wire N__54306;
    wire N__54305;
    wire N__54304;
    wire N__54297;
    wire N__54296;
    wire N__54295;
    wire N__54278;
    wire N__54275;
    wire N__54274;
    wire N__54269;
    wire N__54266;
    wire N__54263;
    wire N__54262;
    wire N__54261;
    wire N__54260;
    wire N__54259;
    wire N__54252;
    wire N__54249;
    wire N__54248;
    wire N__54247;
    wire N__54246;
    wire N__54243;
    wire N__54240;
    wire N__54237;
    wire N__54232;
    wire N__54229;
    wire N__54222;
    wire N__54217;
    wire N__54214;
    wire N__54211;
    wire N__54208;
    wire N__54205;
    wire N__54202;
    wire N__54199;
    wire N__54194;
    wire N__54191;
    wire N__54190;
    wire N__54187;
    wire N__54184;
    wire N__54179;
    wire N__54178;
    wire N__54177;
    wire N__54170;
    wire N__54167;
    wire N__54166;
    wire N__54165;
    wire N__54164;
    wire N__54161;
    wire N__54158;
    wire N__54155;
    wire N__54152;
    wire N__54147;
    wire N__54144;
    wire N__54141;
    wire N__54138;
    wire N__54133;
    wire N__54130;
    wire N__54127;
    wire N__54124;
    wire N__54121;
    wire N__54116;
    wire N__54115;
    wire N__54114;
    wire N__54111;
    wire N__54108;
    wire N__54105;
    wire N__54098;
    wire N__54095;
    wire N__54092;
    wire N__54091;
    wire N__54090;
    wire N__54089;
    wire N__54088;
    wire N__54087;
    wire N__54086;
    wire N__54085;
    wire N__54080;
    wire N__54073;
    wire N__54068;
    wire N__54067;
    wire N__54064;
    wire N__54063;
    wire N__54056;
    wire N__54053;
    wire N__54050;
    wire N__54047;
    wire N__54042;
    wire N__54037;
    wire N__54034;
    wire N__54031;
    wire N__54028;
    wire N__54025;
    wire N__54022;
    wire N__54019;
    wire N__54014;
    wire N__54011;
    wire N__54010;
    wire N__54007;
    wire N__54004;
    wire N__53999;
    wire N__53996;
    wire N__53995;
    wire N__53994;
    wire N__53993;
    wire N__53992;
    wire N__53989;
    wire N__53986;
    wire N__53983;
    wire N__53982;
    wire N__53979;
    wire N__53976;
    wire N__53973;
    wire N__53966;
    wire N__53965;
    wire N__53960;
    wire N__53957;
    wire N__53954;
    wire N__53951;
    wire N__53948;
    wire N__53943;
    wire N__53940;
    wire N__53937;
    wire N__53934;
    wire N__53931;
    wire N__53928;
    wire N__53925;
    wire N__53922;
    wire N__53915;
    wire N__53912;
    wire N__53911;
    wire N__53908;
    wire N__53905;
    wire N__53900;
    wire N__53897;
    wire N__53894;
    wire N__53891;
    wire N__53890;
    wire N__53887;
    wire N__53884;
    wire N__53881;
    wire N__53878;
    wire N__53875;
    wire N__53872;
    wire N__53869;
    wire N__53864;
    wire N__53861;
    wire N__53858;
    wire N__53855;
    wire N__53854;
    wire N__53853;
    wire N__53852;
    wire N__53851;
    wire N__53850;
    wire N__53849;
    wire N__53848;
    wire N__53847;
    wire N__53846;
    wire N__53845;
    wire N__53844;
    wire N__53843;
    wire N__53842;
    wire N__53841;
    wire N__53840;
    wire N__53839;
    wire N__53838;
    wire N__53837;
    wire N__53836;
    wire N__53835;
    wire N__53834;
    wire N__53833;
    wire N__53832;
    wire N__53831;
    wire N__53830;
    wire N__53829;
    wire N__53828;
    wire N__53827;
    wire N__53826;
    wire N__53825;
    wire N__53824;
    wire N__53823;
    wire N__53822;
    wire N__53821;
    wire N__53820;
    wire N__53819;
    wire N__53818;
    wire N__53817;
    wire N__53816;
    wire N__53815;
    wire N__53814;
    wire N__53813;
    wire N__53812;
    wire N__53811;
    wire N__53810;
    wire N__53809;
    wire N__53808;
    wire N__53807;
    wire N__53806;
    wire N__53805;
    wire N__53804;
    wire N__53803;
    wire N__53802;
    wire N__53801;
    wire N__53800;
    wire N__53799;
    wire N__53798;
    wire N__53797;
    wire N__53796;
    wire N__53795;
    wire N__53794;
    wire N__53793;
    wire N__53792;
    wire N__53791;
    wire N__53790;
    wire N__53789;
    wire N__53788;
    wire N__53787;
    wire N__53786;
    wire N__53785;
    wire N__53784;
    wire N__53783;
    wire N__53782;
    wire N__53781;
    wire N__53780;
    wire N__53779;
    wire N__53778;
    wire N__53777;
    wire N__53776;
    wire N__53775;
    wire N__53774;
    wire N__53773;
    wire N__53772;
    wire N__53771;
    wire N__53770;
    wire N__53769;
    wire N__53768;
    wire N__53767;
    wire N__53766;
    wire N__53765;
    wire N__53764;
    wire N__53763;
    wire N__53762;
    wire N__53761;
    wire N__53760;
    wire N__53759;
    wire N__53758;
    wire N__53757;
    wire N__53756;
    wire N__53755;
    wire N__53754;
    wire N__53753;
    wire N__53752;
    wire N__53751;
    wire N__53750;
    wire N__53749;
    wire N__53748;
    wire N__53747;
    wire N__53746;
    wire N__53745;
    wire N__53744;
    wire N__53743;
    wire N__53742;
    wire N__53741;
    wire N__53740;
    wire N__53739;
    wire N__53738;
    wire N__53737;
    wire N__53736;
    wire N__53735;
    wire N__53734;
    wire N__53733;
    wire N__53732;
    wire N__53731;
    wire N__53730;
    wire N__53729;
    wire N__53728;
    wire N__53727;
    wire N__53468;
    wire N__53465;
    wire N__53464;
    wire N__53463;
    wire N__53462;
    wire N__53461;
    wire N__53460;
    wire N__53459;
    wire N__53458;
    wire N__53455;
    wire N__53452;
    wire N__53449;
    wire N__53446;
    wire N__53443;
    wire N__53440;
    wire N__53437;
    wire N__53434;
    wire N__53431;
    wire N__53428;
    wire N__53425;
    wire N__53424;
    wire N__53423;
    wire N__53422;
    wire N__53419;
    wire N__53418;
    wire N__53417;
    wire N__53416;
    wire N__53415;
    wire N__53414;
    wire N__53413;
    wire N__53412;
    wire N__53411;
    wire N__53410;
    wire N__53409;
    wire N__53408;
    wire N__53407;
    wire N__53406;
    wire N__53405;
    wire N__53404;
    wire N__53403;
    wire N__53402;
    wire N__53401;
    wire N__53400;
    wire N__53397;
    wire N__53396;
    wire N__53395;
    wire N__53394;
    wire N__53393;
    wire N__53392;
    wire N__53391;
    wire N__53390;
    wire N__53389;
    wire N__53388;
    wire N__53387;
    wire N__53386;
    wire N__53385;
    wire N__53384;
    wire N__53383;
    wire N__53382;
    wire N__53381;
    wire N__53380;
    wire N__53379;
    wire N__53378;
    wire N__53377;
    wire N__53376;
    wire N__53375;
    wire N__53374;
    wire N__53373;
    wire N__53372;
    wire N__53371;
    wire N__53370;
    wire N__53369;
    wire N__53368;
    wire N__53367;
    wire N__53366;
    wire N__53365;
    wire N__53364;
    wire N__53363;
    wire N__53362;
    wire N__53359;
    wire N__53358;
    wire N__53357;
    wire N__53356;
    wire N__53355;
    wire N__53354;
    wire N__53351;
    wire N__53350;
    wire N__53349;
    wire N__53348;
    wire N__53347;
    wire N__53346;
    wire N__53345;
    wire N__53344;
    wire N__53343;
    wire N__53342;
    wire N__53341;
    wire N__53340;
    wire N__53339;
    wire N__53338;
    wire N__53337;
    wire N__53336;
    wire N__53335;
    wire N__53332;
    wire N__53331;
    wire N__53330;
    wire N__53329;
    wire N__53328;
    wire N__53327;
    wire N__53326;
    wire N__53325;
    wire N__53324;
    wire N__53323;
    wire N__53322;
    wire N__53321;
    wire N__53320;
    wire N__53319;
    wire N__53318;
    wire N__53317;
    wire N__53316;
    wire N__53315;
    wire N__53314;
    wire N__53313;
    wire N__53312;
    wire N__53099;
    wire N__53096;
    wire N__53093;
    wire N__53092;
    wire N__53091;
    wire N__53086;
    wire N__53083;
    wire N__53080;
    wire N__53077;
    wire N__53074;
    wire N__53071;
    wire N__53068;
    wire N__53063;
    wire N__53060;
    wire N__53057;
    wire N__53056;
    wire N__53053;
    wire N__53050;
    wire N__53047;
    wire N__53044;
    wire N__53043;
    wire N__53040;
    wire N__53037;
    wire N__53034;
    wire N__53031;
    wire N__53026;
    wire N__53023;
    wire N__53020;
    wire N__53017;
    wire N__53014;
    wire N__53009;
    wire N__53006;
    wire N__53003;
    wire N__53002;
    wire N__52999;
    wire N__52996;
    wire N__52993;
    wire N__52990;
    wire N__52989;
    wire N__52984;
    wire N__52981;
    wire N__52976;
    wire N__52973;
    wire N__52970;
    wire N__52967;
    wire N__52964;
    wire N__52961;
    wire N__52958;
    wire N__52955;
    wire N__52952;
    wire N__52949;
    wire N__52946;
    wire N__52943;
    wire N__52940;
    wire N__52937;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52925;
    wire N__52922;
    wire N__52919;
    wire N__52916;
    wire N__52913;
    wire N__52910;
    wire N__52907;
    wire N__52904;
    wire N__52901;
    wire N__52898;
    wire N__52895;
    wire N__52892;
    wire N__52889;
    wire N__52886;
    wire N__52883;
    wire N__52880;
    wire N__52877;
    wire N__52874;
    wire N__52871;
    wire N__52868;
    wire N__52865;
    wire N__52862;
    wire N__52859;
    wire N__52856;
    wire N__52853;
    wire N__52850;
    wire N__52847;
    wire N__52844;
    wire N__52841;
    wire N__52838;
    wire N__52835;
    wire N__52832;
    wire N__52831;
    wire N__52830;
    wire N__52827;
    wire N__52824;
    wire N__52821;
    wire N__52814;
    wire N__52811;
    wire N__52808;
    wire N__52805;
    wire N__52802;
    wire N__52799;
    wire N__52796;
    wire N__52795;
    wire N__52794;
    wire N__52793;
    wire N__52792;
    wire N__52791;
    wire N__52790;
    wire N__52789;
    wire N__52788;
    wire N__52787;
    wire N__52786;
    wire N__52785;
    wire N__52784;
    wire N__52783;
    wire N__52782;
    wire N__52781;
    wire N__52764;
    wire N__52747;
    wire N__52742;
    wire N__52739;
    wire N__52738;
    wire N__52737;
    wire N__52736;
    wire N__52735;
    wire N__52734;
    wire N__52731;
    wire N__52726;
    wire N__52719;
    wire N__52716;
    wire N__52711;
    wire N__52708;
    wire N__52703;
    wire N__52700;
    wire N__52699;
    wire N__52698;
    wire N__52695;
    wire N__52690;
    wire N__52687;
    wire N__52684;
    wire N__52681;
    wire N__52678;
    wire N__52675;
    wire N__52672;
    wire N__52667;
    wire N__52664;
    wire N__52661;
    wire N__52658;
    wire N__52655;
    wire N__52652;
    wire N__52649;
    wire N__52648;
    wire N__52643;
    wire N__52640;
    wire N__52637;
    wire N__52634;
    wire N__52631;
    wire N__52628;
    wire N__52625;
    wire N__52622;
    wire N__52621;
    wire N__52618;
    wire N__52615;
    wire N__52612;
    wire N__52609;
    wire N__52606;
    wire N__52601;
    wire N__52600;
    wire N__52597;
    wire N__52594;
    wire N__52591;
    wire N__52588;
    wire N__52585;
    wire N__52580;
    wire N__52579;
    wire N__52576;
    wire N__52573;
    wire N__52570;
    wire N__52567;
    wire N__52564;
    wire N__52559;
    wire N__52558;
    wire N__52555;
    wire N__52550;
    wire N__52547;
    wire N__52544;
    wire N__52543;
    wire N__52538;
    wire N__52535;
    wire N__52532;
    wire N__52531;
    wire N__52526;
    wire N__52523;
    wire N__52520;
    wire N__52519;
    wire N__52514;
    wire N__52511;
    wire N__52508;
    wire N__52505;
    wire N__52504;
    wire N__52501;
    wire N__52498;
    wire N__52495;
    wire N__52490;
    wire N__52487;
    wire N__52484;
    wire N__52481;
    wire N__52478;
    wire N__52475;
    wire N__52472;
    wire N__52469;
    wire N__52466;
    wire N__52463;
    wire N__52462;
    wire N__52459;
    wire N__52456;
    wire N__52455;
    wire N__52454;
    wire N__52451;
    wire N__52448;
    wire N__52445;
    wire N__52442;
    wire N__52439;
    wire N__52432;
    wire N__52427;
    wire N__52426;
    wire N__52425;
    wire N__52424;
    wire N__52423;
    wire N__52422;
    wire N__52421;
    wire N__52420;
    wire N__52419;
    wire N__52418;
    wire N__52417;
    wire N__52416;
    wire N__52413;
    wire N__52408;
    wire N__52405;
    wire N__52402;
    wire N__52401;
    wire N__52400;
    wire N__52397;
    wire N__52394;
    wire N__52389;
    wire N__52388;
    wire N__52387;
    wire N__52384;
    wire N__52379;
    wire N__52376;
    wire N__52375;
    wire N__52374;
    wire N__52373;
    wire N__52372;
    wire N__52371;
    wire N__52370;
    wire N__52369;
    wire N__52368;
    wire N__52367;
    wire N__52366;
    wire N__52365;
    wire N__52364;
    wire N__52363;
    wire N__52362;
    wire N__52361;
    wire N__52358;
    wire N__52355;
    wire N__52352;
    wire N__52347;
    wire N__52344;
    wire N__52339;
    wire N__52332;
    wire N__52329;
    wire N__52326;
    wire N__52323;
    wire N__52320;
    wire N__52307;
    wire N__52304;
    wire N__52291;
    wire N__52284;
    wire N__52275;
    wire N__52268;
    wire N__52253;
    wire N__52250;
    wire N__52247;
    wire N__52244;
    wire N__52241;
    wire N__52240;
    wire N__52239;
    wire N__52238;
    wire N__52237;
    wire N__52236;
    wire N__52235;
    wire N__52234;
    wire N__52233;
    wire N__52230;
    wire N__52227;
    wire N__52224;
    wire N__52223;
    wire N__52222;
    wire N__52221;
    wire N__52216;
    wire N__52215;
    wire N__52214;
    wire N__52213;
    wire N__52212;
    wire N__52211;
    wire N__52210;
    wire N__52209;
    wire N__52208;
    wire N__52207;
    wire N__52206;
    wire N__52205;
    wire N__52204;
    wire N__52201;
    wire N__52198;
    wire N__52197;
    wire N__52196;
    wire N__52191;
    wire N__52190;
    wire N__52189;
    wire N__52188;
    wire N__52187;
    wire N__52184;
    wire N__52181;
    wire N__52178;
    wire N__52173;
    wire N__52170;
    wire N__52167;
    wire N__52154;
    wire N__52141;
    wire N__52136;
    wire N__52131;
    wire N__52128;
    wire N__52125;
    wire N__52122;
    wire N__52117;
    wire N__52112;
    wire N__52109;
    wire N__52106;
    wire N__52095;
    wire N__52090;
    wire N__52073;
    wire N__52072;
    wire N__52069;
    wire N__52068;
    wire N__52065;
    wire N__52062;
    wire N__52059;
    wire N__52058;
    wire N__52055;
    wire N__52050;
    wire N__52047;
    wire N__52044;
    wire N__52039;
    wire N__52036;
    wire N__52033;
    wire N__52030;
    wire N__52027;
    wire N__52022;
    wire N__52021;
    wire N__52016;
    wire N__52013;
    wire N__52010;
    wire N__52009;
    wire N__52006;
    wire N__52003;
    wire N__52000;
    wire N__51995;
    wire N__51992;
    wire N__51989;
    wire N__51986;
    wire N__51985;
    wire N__51980;
    wire N__51977;
    wire N__51974;
    wire N__51973;
    wire N__51968;
    wire N__51965;
    wire N__51962;
    wire N__51959;
    wire N__51956;
    wire N__51953;
    wire N__51950;
    wire N__51949;
    wire N__51946;
    wire N__51943;
    wire N__51938;
    wire N__51935;
    wire N__51932;
    wire N__51929;
    wire N__51928;
    wire N__51925;
    wire N__51922;
    wire N__51919;
    wire N__51916;
    wire N__51911;
    wire N__51908;
    wire N__51907;
    wire N__51902;
    wire N__51899;
    wire N__51896;
    wire N__51895;
    wire N__51890;
    wire N__51887;
    wire N__51884;
    wire N__51881;
    wire N__51878;
    wire N__51877;
    wire N__51874;
    wire N__51871;
    wire N__51866;
    wire N__51863;
    wire N__51860;
    wire N__51859;
    wire N__51856;
    wire N__51853;
    wire N__51850;
    wire N__51847;
    wire N__51842;
    wire N__51841;
    wire N__51836;
    wire N__51833;
    wire N__51830;
    wire N__51829;
    wire N__51824;
    wire N__51821;
    wire N__51818;
    wire N__51815;
    wire N__51814;
    wire N__51813;
    wire N__51810;
    wire N__51805;
    wire N__51804;
    wire N__51801;
    wire N__51798;
    wire N__51795;
    wire N__51790;
    wire N__51785;
    wire N__51782;
    wire N__51781;
    wire N__51780;
    wire N__51777;
    wire N__51772;
    wire N__51771;
    wire N__51768;
    wire N__51765;
    wire N__51762;
    wire N__51757;
    wire N__51752;
    wire N__51749;
    wire N__51748;
    wire N__51747;
    wire N__51746;
    wire N__51743;
    wire N__51740;
    wire N__51737;
    wire N__51734;
    wire N__51731;
    wire N__51728;
    wire N__51723;
    wire N__51720;
    wire N__51717;
    wire N__51714;
    wire N__51707;
    wire N__51706;
    wire N__51705;
    wire N__51702;
    wire N__51699;
    wire N__51696;
    wire N__51693;
    wire N__51690;
    wire N__51689;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51675;
    wire N__51668;
    wire N__51665;
    wire N__51664;
    wire N__51661;
    wire N__51660;
    wire N__51657;
    wire N__51656;
    wire N__51653;
    wire N__51650;
    wire N__51647;
    wire N__51644;
    wire N__51641;
    wire N__51638;
    wire N__51629;
    wire N__51628;
    wire N__51623;
    wire N__51622;
    wire N__51619;
    wire N__51618;
    wire N__51615;
    wire N__51612;
    wire N__51609;
    wire N__51602;
    wire N__51599;
    wire N__51596;
    wire N__51595;
    wire N__51594;
    wire N__51593;
    wire N__51590;
    wire N__51587;
    wire N__51582;
    wire N__51579;
    wire N__51576;
    wire N__51569;
    wire N__51566;
    wire N__51563;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51555;
    wire N__51552;
    wire N__51549;
    wire N__51546;
    wire N__51539;
    wire N__51536;
    wire N__51535;
    wire N__51534;
    wire N__51531;
    wire N__51528;
    wire N__51525;
    wire N__51522;
    wire N__51519;
    wire N__51518;
    wire N__51515;
    wire N__51510;
    wire N__51507;
    wire N__51500;
    wire N__51497;
    wire N__51496;
    wire N__51495;
    wire N__51492;
    wire N__51489;
    wire N__51486;
    wire N__51483;
    wire N__51478;
    wire N__51475;
    wire N__51474;
    wire N__51471;
    wire N__51468;
    wire N__51465;
    wire N__51458;
    wire N__51455;
    wire N__51452;
    wire N__51449;
    wire N__51446;
    wire N__51443;
    wire N__51440;
    wire N__51437;
    wire N__51436;
    wire N__51433;
    wire N__51432;
    wire N__51431;
    wire N__51428;
    wire N__51425;
    wire N__51422;
    wire N__51419;
    wire N__51416;
    wire N__51407;
    wire N__51404;
    wire N__51401;
    wire N__51398;
    wire N__51395;
    wire N__51392;
    wire N__51389;
    wire N__51386;
    wire N__51383;
    wire N__51380;
    wire N__51379;
    wire N__51378;
    wire N__51377;
    wire N__51374;
    wire N__51371;
    wire N__51368;
    wire N__51365;
    wire N__51362;
    wire N__51359;
    wire N__51356;
    wire N__51353;
    wire N__51346;
    wire N__51341;
    wire N__51338;
    wire N__51335;
    wire N__51332;
    wire N__51331;
    wire N__51328;
    wire N__51325;
    wire N__51324;
    wire N__51321;
    wire N__51316;
    wire N__51315;
    wire N__51312;
    wire N__51309;
    wire N__51306;
    wire N__51301;
    wire N__51298;
    wire N__51293;
    wire N__51290;
    wire N__51287;
    wire N__51284;
    wire N__51281;
    wire N__51280;
    wire N__51277;
    wire N__51276;
    wire N__51275;
    wire N__51272;
    wire N__51269;
    wire N__51264;
    wire N__51261;
    wire N__51254;
    wire N__51251;
    wire N__51248;
    wire N__51245;
    wire N__51242;
    wire N__51239;
    wire N__51236;
    wire N__51233;
    wire N__51232;
    wire N__51231;
    wire N__51230;
    wire N__51227;
    wire N__51224;
    wire N__51219;
    wire N__51212;
    wire N__51209;
    wire N__51206;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51196;
    wire N__51193;
    wire N__51190;
    wire N__51189;
    wire N__51188;
    wire N__51185;
    wire N__51182;
    wire N__51179;
    wire N__51176;
    wire N__51167;
    wire N__51164;
    wire N__51161;
    wire N__51158;
    wire N__51155;
    wire N__51152;
    wire N__51149;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51141;
    wire N__51140;
    wire N__51137;
    wire N__51134;
    wire N__51131;
    wire N__51128;
    wire N__51119;
    wire N__51116;
    wire N__51113;
    wire N__51110;
    wire N__51107;
    wire N__51104;
    wire N__51101;
    wire N__51100;
    wire N__51097;
    wire N__51096;
    wire N__51093;
    wire N__51092;
    wire N__51089;
    wire N__51086;
    wire N__51081;
    wire N__51074;
    wire N__51071;
    wire N__51070;
    wire N__51067;
    wire N__51064;
    wire N__51063;
    wire N__51062;
    wire N__51059;
    wire N__51056;
    wire N__51053;
    wire N__51050;
    wire N__51041;
    wire N__51038;
    wire N__51035;
    wire N__51032;
    wire N__51029;
    wire N__51026;
    wire N__51023;
    wire N__51020;
    wire N__51017;
    wire N__51014;
    wire N__51011;
    wire N__51008;
    wire N__51005;
    wire N__51002;
    wire N__50999;
    wire N__50996;
    wire N__50993;
    wire N__50990;
    wire N__50987;
    wire N__50984;
    wire N__50981;
    wire N__50978;
    wire N__50975;
    wire N__50972;
    wire N__50969;
    wire N__50966;
    wire N__50963;
    wire N__50960;
    wire N__50957;
    wire N__50954;
    wire N__50951;
    wire N__50950;
    wire N__50949;
    wire N__50946;
    wire N__50945;
    wire N__50940;
    wire N__50937;
    wire N__50934;
    wire N__50931;
    wire N__50924;
    wire N__50921;
    wire N__50918;
    wire N__50915;
    wire N__50912;
    wire N__50909;
    wire N__50906;
    wire N__50905;
    wire N__50904;
    wire N__50903;
    wire N__50900;
    wire N__50897;
    wire N__50892;
    wire N__50889;
    wire N__50884;
    wire N__50879;
    wire N__50876;
    wire N__50873;
    wire N__50870;
    wire N__50867;
    wire N__50864;
    wire N__50861;
    wire N__50858;
    wire N__50855;
    wire N__50852;
    wire N__50849;
    wire N__50848;
    wire N__50845;
    wire N__50844;
    wire N__50841;
    wire N__50840;
    wire N__50837;
    wire N__50834;
    wire N__50829;
    wire N__50826;
    wire N__50823;
    wire N__50820;
    wire N__50813;
    wire N__50810;
    wire N__50807;
    wire N__50804;
    wire N__50801;
    wire N__50798;
    wire N__50795;
    wire N__50794;
    wire N__50793;
    wire N__50790;
    wire N__50787;
    wire N__50786;
    wire N__50783;
    wire N__50780;
    wire N__50777;
    wire N__50772;
    wire N__50765;
    wire N__50762;
    wire N__50759;
    wire N__50756;
    wire N__50753;
    wire N__50750;
    wire N__50749;
    wire N__50748;
    wire N__50747;
    wire N__50744;
    wire N__50741;
    wire N__50736;
    wire N__50731;
    wire N__50728;
    wire N__50725;
    wire N__50720;
    wire N__50717;
    wire N__50714;
    wire N__50711;
    wire N__50708;
    wire N__50705;
    wire N__50702;
    wire N__50699;
    wire N__50696;
    wire N__50693;
    wire N__50692;
    wire N__50689;
    wire N__50686;
    wire N__50685;
    wire N__50682;
    wire N__50681;
    wire N__50678;
    wire N__50675;
    wire N__50672;
    wire N__50669;
    wire N__50664;
    wire N__50661;
    wire N__50658;
    wire N__50655;
    wire N__50648;
    wire N__50645;
    wire N__50642;
    wire N__50639;
    wire N__50636;
    wire N__50633;
    wire N__50630;
    wire N__50629;
    wire N__50626;
    wire N__50623;
    wire N__50622;
    wire N__50619;
    wire N__50618;
    wire N__50615;
    wire N__50612;
    wire N__50609;
    wire N__50606;
    wire N__50603;
    wire N__50594;
    wire N__50591;
    wire N__50588;
    wire N__50585;
    wire N__50582;
    wire N__50579;
    wire N__50578;
    wire N__50575;
    wire N__50572;
    wire N__50571;
    wire N__50570;
    wire N__50565;
    wire N__50562;
    wire N__50559;
    wire N__50556;
    wire N__50549;
    wire N__50546;
    wire N__50543;
    wire N__50540;
    wire N__50537;
    wire N__50534;
    wire N__50531;
    wire N__50528;
    wire N__50527;
    wire N__50526;
    wire N__50523;
    wire N__50522;
    wire N__50517;
    wire N__50514;
    wire N__50511;
    wire N__50508;
    wire N__50501;
    wire N__50498;
    wire N__50495;
    wire N__50492;
    wire N__50489;
    wire N__50486;
    wire N__50483;
    wire N__50480;
    wire N__50477;
    wire N__50474;
    wire N__50471;
    wire N__50468;
    wire N__50465;
    wire N__50462;
    wire N__50459;
    wire N__50456;
    wire N__50453;
    wire N__50450;
    wire N__50447;
    wire N__50444;
    wire N__50441;
    wire N__50438;
    wire N__50435;
    wire N__50432;
    wire N__50429;
    wire N__50426;
    wire N__50423;
    wire N__50420;
    wire N__50417;
    wire N__50414;
    wire N__50411;
    wire N__50408;
    wire N__50405;
    wire N__50402;
    wire N__50399;
    wire N__50396;
    wire N__50393;
    wire N__50390;
    wire N__50387;
    wire N__50384;
    wire N__50381;
    wire N__50378;
    wire N__50375;
    wire N__50374;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50360;
    wire N__50357;
    wire N__50354;
    wire N__50353;
    wire N__50350;
    wire N__50347;
    wire N__50344;
    wire N__50339;
    wire N__50336;
    wire N__50333;
    wire N__50330;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50320;
    wire N__50315;
    wire N__50312;
    wire N__50309;
    wire N__50306;
    wire N__50303;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50282;
    wire N__50279;
    wire N__50278;
    wire N__50275;
    wire N__50272;
    wire N__50269;
    wire N__50264;
    wire N__50261;
    wire N__50258;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50237;
    wire N__50234;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50219;
    wire N__50216;
    wire N__50213;
    wire N__50210;
    wire N__50207;
    wire N__50206;
    wire N__50203;
    wire N__50200;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50186;
    wire N__50185;
    wire N__50182;
    wire N__50179;
    wire N__50176;
    wire N__50171;
    wire N__50168;
    wire N__50165;
    wire N__50164;
    wire N__50159;
    wire N__50158;
    wire N__50155;
    wire N__50152;
    wire N__50149;
    wire N__50146;
    wire N__50141;
    wire N__50138;
    wire N__50137;
    wire N__50136;
    wire N__50135;
    wire N__50132;
    wire N__50127;
    wire N__50126;
    wire N__50125;
    wire N__50122;
    wire N__50121;
    wire N__50120;
    wire N__50119;
    wire N__50118;
    wire N__50117;
    wire N__50112;
    wire N__50111;
    wire N__50108;
    wire N__50107;
    wire N__50106;
    wire N__50105;
    wire N__50104;
    wire N__50103;
    wire N__50102;
    wire N__50101;
    wire N__50100;
    wire N__50099;
    wire N__50098;
    wire N__50097;
    wire N__50096;
    wire N__50095;
    wire N__50092;
    wire N__50091;
    wire N__50090;
    wire N__50089;
    wire N__50088;
    wire N__50087;
    wire N__50086;
    wire N__50085;
    wire N__50084;
    wire N__50083;
    wire N__50082;
    wire N__50081;
    wire N__50068;
    wire N__50065;
    wire N__50060;
    wire N__50059;
    wire N__50050;
    wire N__50049;
    wire N__50046;
    wire N__50033;
    wire N__50028;
    wire N__50025;
    wire N__50022;
    wire N__50021;
    wire N__50004;
    wire N__49999;
    wire N__49998;
    wire N__49997;
    wire N__49996;
    wire N__49995;
    wire N__49994;
    wire N__49993;
    wire N__49992;
    wire N__49991;
    wire N__49990;
    wire N__49989;
    wire N__49988;
    wire N__49987;
    wire N__49986;
    wire N__49985;
    wire N__49982;
    wire N__49981;
    wire N__49980;
    wire N__49979;
    wire N__49978;
    wire N__49973;
    wire N__49970;
    wire N__49967;
    wire N__49964;
    wire N__49959;
    wire N__49952;
    wire N__49951;
    wire N__49950;
    wire N__49949;
    wire N__49948;
    wire N__49947;
    wire N__49946;
    wire N__49945;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49941;
    wire N__49940;
    wire N__49937;
    wire N__49936;
    wire N__49935;
    wire N__49930;
    wire N__49923;
    wire N__49912;
    wire N__49899;
    wire N__49896;
    wire N__49887;
    wire N__49884;
    wire N__49881;
    wire N__49878;
    wire N__49871;
    wire N__49854;
    wire N__49851;
    wire N__49838;
    wire N__49835;
    wire N__49824;
    wire N__49805;
    wire N__49804;
    wire N__49801;
    wire N__49796;
    wire N__49793;
    wire N__49792;
    wire N__49789;
    wire N__49786;
    wire N__49785;
    wire N__49782;
    wire N__49779;
    wire N__49776;
    wire N__49769;
    wire N__49768;
    wire N__49767;
    wire N__49766;
    wire N__49765;
    wire N__49762;
    wire N__49761;
    wire N__49760;
    wire N__49759;
    wire N__49758;
    wire N__49757;
    wire N__49756;
    wire N__49753;
    wire N__49752;
    wire N__49751;
    wire N__49750;
    wire N__49747;
    wire N__49746;
    wire N__49743;
    wire N__49740;
    wire N__49737;
    wire N__49736;
    wire N__49733;
    wire N__49730;
    wire N__49729;
    wire N__49728;
    wire N__49727;
    wire N__49724;
    wire N__49723;
    wire N__49720;
    wire N__49719;
    wire N__49718;
    wire N__49717;
    wire N__49716;
    wire N__49715;
    wire N__49714;
    wire N__49713;
    wire N__49712;
    wire N__49709;
    wire N__49708;
    wire N__49707;
    wire N__49706;
    wire N__49705;
    wire N__49702;
    wire N__49685;
    wire N__49682;
    wire N__49667;
    wire N__49662;
    wire N__49651;
    wire N__49650;
    wire N__49649;
    wire N__49640;
    wire N__49639;
    wire N__49636;
    wire N__49635;
    wire N__49634;
    wire N__49631;
    wire N__49628;
    wire N__49625;
    wire N__49624;
    wire N__49623;
    wire N__49622;
    wire N__49621;
    wire N__49620;
    wire N__49619;
    wire N__49618;
    wire N__49617;
    wire N__49616;
    wire N__49615;
    wire N__49614;
    wire N__49613;
    wire N__49612;
    wire N__49609;
    wire N__49606;
    wire N__49597;
    wire N__49592;
    wire N__49589;
    wire N__49586;
    wire N__49583;
    wire N__49572;
    wire N__49569;
    wire N__49564;
    wire N__49563;
    wire N__49562;
    wire N__49561;
    wire N__49560;
    wire N__49559;
    wire N__49558;
    wire N__49557;
    wire N__49556;
    wire N__49555;
    wire N__49554;
    wire N__49553;
    wire N__49552;
    wire N__49551;
    wire N__49550;
    wire N__49549;
    wire N__49548;
    wire N__49547;
    wire N__49546;
    wire N__49545;
    wire N__49544;
    wire N__49543;
    wire N__49542;
    wire N__49541;
    wire N__49540;
    wire N__49539;
    wire N__49538;
    wire N__49535;
    wire N__49534;
    wire N__49531;
    wire N__49530;
    wire N__49527;
    wire N__49526;
    wire N__49523;
    wire N__49522;
    wire N__49519;
    wire N__49518;
    wire N__49515;
    wire N__49514;
    wire N__49511;
    wire N__49510;
    wire N__49509;
    wire N__49508;
    wire N__49507;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49503;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49499;
    wire N__49496;
    wire N__49495;
    wire N__49492;
    wire N__49491;
    wire N__49488;
    wire N__49487;
    wire N__49484;
    wire N__49477;
    wire N__49468;
    wire N__49463;
    wire N__49460;
    wire N__49459;
    wire N__49456;
    wire N__49441;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49429;
    wire N__49428;
    wire N__49425;
    wire N__49424;
    wire N__49421;
    wire N__49420;
    wire N__49417;
    wire N__49416;
    wire N__49413;
    wire N__49412;
    wire N__49409;
    wire N__49408;
    wire N__49405;
    wire N__49404;
    wire N__49399;
    wire N__49390;
    wire N__49375;
    wire N__49358;
    wire N__49355;
    wire N__49354;
    wire N__49351;
    wire N__49350;
    wire N__49347;
    wire N__49346;
    wire N__49343;
    wire N__49342;
    wire N__49339;
    wire N__49338;
    wire N__49335;
    wire N__49334;
    wire N__49331;
    wire N__49330;
    wire N__49327;
    wire N__49326;
    wire N__49323;
    wire N__49322;
    wire N__49319;
    wire N__49318;
    wire N__49315;
    wire N__49314;
    wire N__49301;
    wire N__49298;
    wire N__49295;
    wire N__49292;
    wire N__49287;
    wire N__49282;
    wire N__49277;
    wire N__49260;
    wire N__49243;
    wire N__49234;
    wire N__49217;
    wire N__49200;
    wire N__49187;
    wire N__49184;
    wire N__49157;
    wire N__49154;
    wire N__49151;
    wire N__49148;
    wire N__49145;
    wire N__49144;
    wire N__49143;
    wire N__49138;
    wire N__49135;
    wire N__49130;
    wire N__49129;
    wire N__49128;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49118;
    wire N__49115;
    wire N__49110;
    wire N__49107;
    wire N__49104;
    wire N__49097;
    wire N__49094;
    wire N__49091;
    wire N__49088;
    wire N__49085;
    wire N__49084;
    wire N__49083;
    wire N__49080;
    wire N__49075;
    wire N__49072;
    wire N__49069;
    wire N__49064;
    wire N__49063;
    wire N__49062;
    wire N__49061;
    wire N__49058;
    wire N__49055;
    wire N__49052;
    wire N__49049;
    wire N__49046;
    wire N__49037;
    wire N__49036;
    wire N__49033;
    wire N__49032;
    wire N__49031;
    wire N__49028;
    wire N__49023;
    wire N__49020;
    wire N__49017;
    wire N__49010;
    wire N__49007;
    wire N__49004;
    wire N__49001;
    wire N__48998;
    wire N__48995;
    wire N__48992;
    wire N__48989;
    wire N__48986;
    wire N__48983;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48968;
    wire N__48965;
    wire N__48964;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48950;
    wire N__48947;
    wire N__48944;
    wire N__48941;
    wire N__48940;
    wire N__48937;
    wire N__48934;
    wire N__48931;
    wire N__48926;
    wire N__48923;
    wire N__48920;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48910;
    wire N__48905;
    wire N__48902;
    wire N__48899;
    wire N__48896;
    wire N__48893;
    wire N__48890;
    wire N__48887;
    wire N__48884;
    wire N__48881;
    wire N__48878;
    wire N__48877;
    wire N__48872;
    wire N__48871;
    wire N__48870;
    wire N__48867;
    wire N__48862;
    wire N__48859;
    wire N__48854;
    wire N__48853;
    wire N__48850;
    wire N__48849;
    wire N__48842;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48830;
    wire N__48827;
    wire N__48824;
    wire N__48821;
    wire N__48818;
    wire N__48817;
    wire N__48816;
    wire N__48815;
    wire N__48812;
    wire N__48809;
    wire N__48806;
    wire N__48803;
    wire N__48794;
    wire N__48793;
    wire N__48792;
    wire N__48791;
    wire N__48784;
    wire N__48781;
    wire N__48776;
    wire N__48775;
    wire N__48774;
    wire N__48773;
    wire N__48772;
    wire N__48771;
    wire N__48770;
    wire N__48769;
    wire N__48768;
    wire N__48767;
    wire N__48766;
    wire N__48765;
    wire N__48756;
    wire N__48755;
    wire N__48754;
    wire N__48753;
    wire N__48752;
    wire N__48751;
    wire N__48750;
    wire N__48749;
    wire N__48748;
    wire N__48747;
    wire N__48746;
    wire N__48745;
    wire N__48744;
    wire N__48735;
    wire N__48726;
    wire N__48725;
    wire N__48724;
    wire N__48723;
    wire N__48722;
    wire N__48721;
    wire N__48720;
    wire N__48717;
    wire N__48708;
    wire N__48699;
    wire N__48690;
    wire N__48685;
    wire N__48680;
    wire N__48671;
    wire N__48668;
    wire N__48659;
    wire N__48650;
    wire N__48647;
    wire N__48644;
    wire N__48641;
    wire N__48638;
    wire N__48635;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48623;
    wire N__48620;
    wire N__48617;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48605;
    wire N__48602;
    wire N__48599;
    wire N__48596;
    wire N__48593;
    wire N__48590;
    wire N__48587;
    wire N__48584;
    wire N__48581;
    wire N__48578;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48563;
    wire N__48560;
    wire N__48557;
    wire N__48554;
    wire N__48551;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48539;
    wire N__48536;
    wire N__48533;
    wire N__48530;
    wire N__48527;
    wire N__48524;
    wire N__48521;
    wire N__48518;
    wire N__48515;
    wire N__48512;
    wire N__48509;
    wire N__48506;
    wire N__48503;
    wire N__48500;
    wire N__48497;
    wire N__48494;
    wire N__48491;
    wire N__48488;
    wire N__48485;
    wire N__48482;
    wire N__48479;
    wire N__48476;
    wire N__48473;
    wire N__48470;
    wire N__48467;
    wire N__48464;
    wire N__48461;
    wire N__48458;
    wire N__48455;
    wire N__48452;
    wire N__48449;
    wire N__48446;
    wire N__48443;
    wire N__48440;
    wire N__48437;
    wire N__48434;
    wire N__48431;
    wire N__48428;
    wire N__48425;
    wire N__48422;
    wire N__48419;
    wire N__48416;
    wire N__48413;
    wire N__48410;
    wire N__48407;
    wire N__48404;
    wire N__48401;
    wire N__48398;
    wire N__48395;
    wire N__48392;
    wire N__48389;
    wire N__48386;
    wire N__48383;
    wire N__48380;
    wire N__48377;
    wire N__48374;
    wire N__48371;
    wire N__48368;
    wire N__48365;
    wire N__48362;
    wire N__48359;
    wire N__48356;
    wire N__48353;
    wire N__48350;
    wire N__48347;
    wire N__48344;
    wire N__48341;
    wire N__48338;
    wire N__48335;
    wire N__48332;
    wire N__48329;
    wire N__48326;
    wire N__48323;
    wire N__48320;
    wire N__48317;
    wire N__48314;
    wire N__48311;
    wire N__48308;
    wire N__48305;
    wire N__48302;
    wire N__48299;
    wire N__48296;
    wire N__48293;
    wire N__48290;
    wire N__48287;
    wire N__48284;
    wire N__48281;
    wire N__48278;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48263;
    wire N__48260;
    wire N__48257;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48242;
    wire N__48239;
    wire N__48236;
    wire N__48233;
    wire N__48230;
    wire N__48227;
    wire N__48224;
    wire N__48221;
    wire N__48218;
    wire N__48215;
    wire N__48212;
    wire N__48209;
    wire N__48206;
    wire N__48203;
    wire N__48200;
    wire N__48197;
    wire N__48194;
    wire N__48191;
    wire N__48188;
    wire N__48185;
    wire N__48182;
    wire N__48179;
    wire N__48176;
    wire N__48173;
    wire N__48170;
    wire N__48167;
    wire N__48164;
    wire N__48161;
    wire N__48158;
    wire N__48155;
    wire N__48152;
    wire N__48149;
    wire N__48146;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48128;
    wire N__48125;
    wire N__48122;
    wire N__48119;
    wire N__48116;
    wire N__48113;
    wire N__48110;
    wire N__48107;
    wire N__48104;
    wire N__48101;
    wire N__48098;
    wire N__48095;
    wire N__48092;
    wire N__48089;
    wire N__48086;
    wire N__48083;
    wire N__48080;
    wire N__48077;
    wire N__48074;
    wire N__48071;
    wire N__48068;
    wire N__48065;
    wire N__48062;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48047;
    wire N__48044;
    wire N__48041;
    wire N__48038;
    wire N__48035;
    wire N__48032;
    wire N__48029;
    wire N__48026;
    wire N__48023;
    wire N__48020;
    wire N__48017;
    wire N__48014;
    wire N__48011;
    wire N__48008;
    wire N__48005;
    wire N__48002;
    wire N__47999;
    wire N__47996;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47984;
    wire N__47981;
    wire N__47978;
    wire N__47975;
    wire N__47972;
    wire N__47969;
    wire N__47966;
    wire N__47963;
    wire N__47960;
    wire N__47957;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47945;
    wire N__47942;
    wire N__47939;
    wire N__47936;
    wire N__47933;
    wire N__47930;
    wire N__47927;
    wire N__47924;
    wire N__47921;
    wire N__47918;
    wire N__47915;
    wire N__47912;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47864;
    wire N__47861;
    wire N__47858;
    wire N__47855;
    wire N__47852;
    wire N__47849;
    wire N__47846;
    wire N__47843;
    wire N__47840;
    wire N__47837;
    wire N__47834;
    wire N__47831;
    wire N__47828;
    wire N__47825;
    wire N__47822;
    wire N__47819;
    wire N__47816;
    wire N__47813;
    wire N__47810;
    wire N__47807;
    wire N__47804;
    wire N__47801;
    wire N__47798;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47786;
    wire N__47783;
    wire N__47780;
    wire N__47777;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47723;
    wire N__47720;
    wire N__47717;
    wire N__47714;
    wire N__47711;
    wire N__47708;
    wire N__47705;
    wire N__47702;
    wire N__47699;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47687;
    wire N__47686;
    wire N__47685;
    wire N__47682;
    wire N__47681;
    wire N__47680;
    wire N__47675;
    wire N__47672;
    wire N__47671;
    wire N__47666;
    wire N__47665;
    wire N__47664;
    wire N__47663;
    wire N__47662;
    wire N__47661;
    wire N__47660;
    wire N__47659;
    wire N__47656;
    wire N__47653;
    wire N__47652;
    wire N__47651;
    wire N__47650;
    wire N__47649;
    wire N__47648;
    wire N__47647;
    wire N__47644;
    wire N__47641;
    wire N__47636;
    wire N__47625;
    wire N__47624;
    wire N__47623;
    wire N__47622;
    wire N__47621;
    wire N__47620;
    wire N__47619;
    wire N__47618;
    wire N__47617;
    wire N__47616;
    wire N__47615;
    wire N__47614;
    wire N__47613;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47593;
    wire N__47584;
    wire N__47567;
    wire N__47556;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47525;
    wire N__47522;
    wire N__47519;
    wire N__47516;
    wire N__47513;
    wire N__47510;
    wire N__47507;
    wire N__47504;
    wire N__47501;
    wire N__47498;
    wire N__47495;
    wire N__47492;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47480;
    wire N__47477;
    wire N__47474;
    wire N__47471;
    wire N__47468;
    wire N__47465;
    wire N__47462;
    wire N__47459;
    wire N__47456;
    wire N__47453;
    wire N__47450;
    wire N__47447;
    wire N__47444;
    wire N__47441;
    wire N__47438;
    wire N__47435;
    wire N__47432;
    wire N__47429;
    wire N__47426;
    wire N__47423;
    wire N__47420;
    wire N__47417;
    wire N__47414;
    wire N__47411;
    wire N__47408;
    wire N__47405;
    wire N__47402;
    wire N__47399;
    wire N__47396;
    wire N__47393;
    wire N__47390;
    wire N__47387;
    wire N__47384;
    wire N__47381;
    wire N__47378;
    wire N__47375;
    wire N__47372;
    wire N__47369;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47348;
    wire N__47345;
    wire N__47342;
    wire N__47339;
    wire N__47336;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47324;
    wire N__47321;
    wire N__47318;
    wire N__47315;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47303;
    wire N__47300;
    wire N__47297;
    wire N__47294;
    wire N__47291;
    wire N__47288;
    wire N__47285;
    wire N__47282;
    wire N__47279;
    wire N__47276;
    wire N__47273;
    wire N__47270;
    wire N__47267;
    wire N__47264;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47252;
    wire N__47249;
    wire N__47246;
    wire N__47243;
    wire N__47240;
    wire N__47237;
    wire N__47234;
    wire N__47231;
    wire N__47228;
    wire N__47225;
    wire N__47222;
    wire N__47219;
    wire N__47216;
    wire N__47213;
    wire N__47210;
    wire N__47207;
    wire N__47204;
    wire N__47201;
    wire N__47198;
    wire N__47195;
    wire N__47192;
    wire N__47189;
    wire N__47186;
    wire N__47183;
    wire N__47180;
    wire N__47177;
    wire N__47174;
    wire N__47171;
    wire N__47168;
    wire N__47165;
    wire N__47162;
    wire N__47159;
    wire N__47156;
    wire N__47153;
    wire N__47150;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47135;
    wire N__47132;
    wire N__47129;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47117;
    wire N__47114;
    wire N__47111;
    wire N__47108;
    wire N__47105;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47084;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47054;
    wire N__47051;
    wire N__47048;
    wire N__47045;
    wire N__47042;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47030;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47015;
    wire N__47012;
    wire N__47009;
    wire N__47006;
    wire N__47003;
    wire N__47000;
    wire N__46997;
    wire N__46994;
    wire N__46991;
    wire N__46988;
    wire N__46985;
    wire N__46982;
    wire N__46979;
    wire N__46976;
    wire N__46973;
    wire N__46970;
    wire N__46967;
    wire N__46964;
    wire N__46961;
    wire N__46958;
    wire N__46955;
    wire N__46952;
    wire N__46949;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46937;
    wire N__46934;
    wire N__46931;
    wire N__46928;
    wire N__46925;
    wire N__46922;
    wire N__46919;
    wire N__46916;
    wire N__46913;
    wire N__46910;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46898;
    wire N__46895;
    wire N__46892;
    wire N__46889;
    wire N__46886;
    wire N__46883;
    wire N__46880;
    wire N__46877;
    wire N__46874;
    wire N__46871;
    wire N__46868;
    wire N__46865;
    wire N__46862;
    wire N__46859;
    wire N__46856;
    wire N__46853;
    wire N__46850;
    wire N__46847;
    wire N__46844;
    wire N__46841;
    wire N__46838;
    wire N__46835;
    wire N__46832;
    wire N__46829;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46821;
    wire N__46818;
    wire N__46815;
    wire N__46812;
    wire N__46805;
    wire N__46802;
    wire N__46799;
    wire N__46796;
    wire N__46793;
    wire N__46790;
    wire N__46787;
    wire N__46784;
    wire N__46781;
    wire N__46778;
    wire N__46775;
    wire N__46772;
    wire N__46769;
    wire N__46766;
    wire N__46763;
    wire N__46760;
    wire N__46757;
    wire N__46754;
    wire N__46751;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46739;
    wire N__46736;
    wire N__46733;
    wire N__46730;
    wire N__46727;
    wire N__46724;
    wire N__46721;
    wire N__46718;
    wire N__46715;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46700;
    wire N__46697;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46685;
    wire N__46682;
    wire N__46679;
    wire N__46676;
    wire N__46673;
    wire N__46670;
    wire N__46667;
    wire N__46664;
    wire N__46661;
    wire N__46658;
    wire N__46655;
    wire N__46652;
    wire N__46649;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46619;
    wire N__46616;
    wire N__46613;
    wire N__46610;
    wire N__46607;
    wire N__46604;
    wire N__46601;
    wire N__46598;
    wire N__46595;
    wire N__46592;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46580;
    wire N__46577;
    wire N__46574;
    wire N__46571;
    wire N__46568;
    wire N__46565;
    wire N__46562;
    wire N__46559;
    wire N__46556;
    wire N__46553;
    wire N__46550;
    wire N__46547;
    wire N__46544;
    wire N__46541;
    wire N__46538;
    wire N__46535;
    wire N__46532;
    wire N__46529;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46511;
    wire N__46508;
    wire N__46505;
    wire N__46502;
    wire N__46499;
    wire N__46496;
    wire N__46493;
    wire N__46490;
    wire N__46487;
    wire N__46484;
    wire N__46481;
    wire N__46478;
    wire N__46475;
    wire N__46472;
    wire N__46469;
    wire N__46466;
    wire N__46463;
    wire N__46460;
    wire N__46457;
    wire N__46454;
    wire N__46451;
    wire N__46448;
    wire N__46445;
    wire N__46442;
    wire N__46439;
    wire N__46436;
    wire N__46433;
    wire N__46430;
    wire N__46427;
    wire N__46426;
    wire N__46425;
    wire N__46422;
    wire N__46421;
    wire N__46420;
    wire N__46419;
    wire N__46414;
    wire N__46409;
    wire N__46406;
    wire N__46403;
    wire N__46400;
    wire N__46397;
    wire N__46394;
    wire N__46391;
    wire N__46388;
    wire N__46381;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46367;
    wire N__46364;
    wire N__46361;
    wire N__46358;
    wire N__46355;
    wire N__46352;
    wire N__46349;
    wire N__46346;
    wire N__46343;
    wire N__46340;
    wire N__46337;
    wire N__46334;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46322;
    wire N__46319;
    wire N__46316;
    wire N__46313;
    wire N__46310;
    wire N__46307;
    wire N__46304;
    wire N__46301;
    wire N__46298;
    wire N__46295;
    wire N__46292;
    wire N__46289;
    wire N__46286;
    wire N__46283;
    wire N__46280;
    wire N__46277;
    wire N__46274;
    wire N__46271;
    wire N__46268;
    wire N__46265;
    wire N__46262;
    wire N__46259;
    wire N__46256;
    wire N__46253;
    wire N__46250;
    wire N__46247;
    wire N__46244;
    wire N__46241;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46229;
    wire N__46226;
    wire N__46223;
    wire N__46220;
    wire N__46217;
    wire N__46214;
    wire N__46211;
    wire N__46208;
    wire N__46205;
    wire N__46202;
    wire N__46199;
    wire N__46196;
    wire N__46193;
    wire N__46190;
    wire N__46187;
    wire N__46184;
    wire N__46181;
    wire N__46178;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46136;
    wire N__46133;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46105;
    wire N__46102;
    wire N__46097;
    wire N__46094;
    wire N__46093;
    wire N__46088;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46073;
    wire N__46070;
    wire N__46069;
    wire N__46064;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46049;
    wire N__46046;
    wire N__46043;
    wire N__46040;
    wire N__46037;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46027;
    wire N__46022;
    wire N__46019;
    wire N__46016;
    wire N__46013;
    wire N__46010;
    wire N__46009;
    wire N__46006;
    wire N__46003;
    wire N__46000;
    wire N__45995;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45983;
    wire N__45980;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45970;
    wire N__45967;
    wire N__45962;
    wire N__45959;
    wire N__45956;
    wire N__45953;
    wire N__45950;
    wire N__45947;
    wire N__45944;
    wire N__45943;
    wire N__45940;
    wire N__45935;
    wire N__45932;
    wire N__45931;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45921;
    wire N__45916;
    wire N__45911;
    wire N__45910;
    wire N__45905;
    wire N__45904;
    wire N__45901;
    wire N__45898;
    wire N__45895;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45883;
    wire N__45882;
    wire N__45879;
    wire N__45876;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45862;
    wire N__45859;
    wire N__45854;
    wire N__45851;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45823;
    wire N__45820;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45808;
    wire N__45805;
    wire N__45802;
    wire N__45801;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45785;
    wire N__45782;
    wire N__45781;
    wire N__45776;
    wire N__45775;
    wire N__45772;
    wire N__45769;
    wire N__45766;
    wire N__45761;
    wire N__45758;
    wire N__45755;
    wire N__45754;
    wire N__45751;
    wire N__45748;
    wire N__45747;
    wire N__45742;
    wire N__45739;
    wire N__45736;
    wire N__45731;
    wire N__45728;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45716;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45706;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45694;
    wire N__45691;
    wire N__45688;
    wire N__45687;
    wire N__45682;
    wire N__45679;
    wire N__45676;
    wire N__45671;
    wire N__45668;
    wire N__45667;
    wire N__45662;
    wire N__45661;
    wire N__45658;
    wire N__45655;
    wire N__45652;
    wire N__45647;
    wire N__45644;
    wire N__45643;
    wire N__45638;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45628;
    wire N__45623;
    wire N__45620;
    wire N__45617;
    wire N__45616;
    wire N__45615;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45600;
    wire N__45595;
    wire N__45592;
    wire N__45587;
    wire N__45584;
    wire N__45583;
    wire N__45580;
    wire N__45577;
    wire N__45574;
    wire N__45571;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45548;
    wire N__45545;
    wire N__45542;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45534;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45518;
    wire N__45515;
    wire N__45514;
    wire N__45509;
    wire N__45508;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45494;
    wire N__45491;
    wire N__45490;
    wire N__45485;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45470;
    wire N__45467;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45455;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45440;
    wire N__45437;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45425;
    wire N__45424;
    wire N__45421;
    wire N__45418;
    wire N__45415;
    wire N__45410;
    wire N__45407;
    wire N__45406;
    wire N__45405;
    wire N__45404;
    wire N__45403;
    wire N__45402;
    wire N__45401;
    wire N__45400;
    wire N__45399;
    wire N__45398;
    wire N__45397;
    wire N__45396;
    wire N__45395;
    wire N__45394;
    wire N__45393;
    wire N__45392;
    wire N__45391;
    wire N__45390;
    wire N__45389;
    wire N__45388;
    wire N__45387;
    wire N__45386;
    wire N__45385;
    wire N__45384;
    wire N__45383;
    wire N__45382;
    wire N__45381;
    wire N__45380;
    wire N__45379;
    wire N__45378;
    wire N__45369;
    wire N__45364;
    wire N__45355;
    wire N__45346;
    wire N__45337;
    wire N__45328;
    wire N__45319;
    wire N__45310;
    wire N__45303;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45283;
    wire N__45280;
    wire N__45277;
    wire N__45274;
    wire N__45269;
    wire N__45268;
    wire N__45267;
    wire N__45264;
    wire N__45261;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45251;
    wire N__45248;
    wire N__45243;
    wire N__45240;
    wire N__45233;
    wire N__45230;
    wire N__45227;
    wire N__45224;
    wire N__45223;
    wire N__45220;
    wire N__45217;
    wire N__45216;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45202;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45160;
    wire N__45155;
    wire N__45152;
    wire N__45151;
    wire N__45146;
    wire N__45145;
    wire N__45142;
    wire N__45139;
    wire N__45136;
    wire N__45131;
    wire N__45128;
    wire N__45127;
    wire N__45122;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45112;
    wire N__45107;
    wire N__45104;
    wire N__45103;
    wire N__45100;
    wire N__45097;
    wire N__45092;
    wire N__45091;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45077;
    wire N__45074;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45062;
    wire N__45061;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45040;
    wire N__45037;
    wire N__45034;
    wire N__45033;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45017;
    wire N__45014;
    wire N__45013;
    wire N__45010;
    wire N__45007;
    wire N__45006;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44990;
    wire N__44987;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44979;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44963;
    wire N__44960;
    wire N__44957;
    wire N__44956;
    wire N__44955;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44941;
    wire N__44936;
    wire N__44933;
    wire N__44930;
    wire N__44929;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44914;
    wire N__44909;
    wire N__44906;
    wire N__44903;
    wire N__44900;
    wire N__44899;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44876;
    wire N__44873;
    wire N__44870;
    wire N__44867;
    wire N__44866;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44843;
    wire N__44840;
    wire N__44839;
    wire N__44838;
    wire N__44833;
    wire N__44830;
    wire N__44827;
    wire N__44822;
    wire N__44819;
    wire N__44818;
    wire N__44817;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44801;
    wire N__44798;
    wire N__44795;
    wire N__44794;
    wire N__44791;
    wire N__44788;
    wire N__44785;
    wire N__44780;
    wire N__44777;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44765;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44750;
    wire N__44747;
    wire N__44746;
    wire N__44743;
    wire N__44740;
    wire N__44735;
    wire N__44734;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44720;
    wire N__44717;
    wire N__44714;
    wire N__44713;
    wire N__44710;
    wire N__44707;
    wire N__44706;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44690;
    wire N__44687;
    wire N__44686;
    wire N__44681;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44671;
    wire N__44666;
    wire N__44663;
    wire N__44660;
    wire N__44657;
    wire N__44656;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44643;
    wire N__44640;
    wire N__44633;
    wire N__44630;
    wire N__44627;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44619;
    wire N__44616;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44597;
    wire N__44594;
    wire N__44593;
    wire N__44588;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44573;
    wire N__44570;
    wire N__44569;
    wire N__44564;
    wire N__44563;
    wire N__44560;
    wire N__44557;
    wire N__44554;
    wire N__44549;
    wire N__44546;
    wire N__44545;
    wire N__44540;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44525;
    wire N__44522;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44510;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44495;
    wire N__44492;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44480;
    wire N__44479;
    wire N__44476;
    wire N__44473;
    wire N__44470;
    wire N__44465;
    wire N__44462;
    wire N__44459;
    wire N__44458;
    wire N__44455;
    wire N__44452;
    wire N__44451;
    wire N__44446;
    wire N__44443;
    wire N__44440;
    wire N__44435;
    wire N__44432;
    wire N__44429;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44421;
    wire N__44416;
    wire N__44413;
    wire N__44410;
    wire N__44405;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44395;
    wire N__44394;
    wire N__44391;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44363;
    wire N__44362;
    wire N__44361;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44347;
    wire N__44342;
    wire N__44339;
    wire N__44338;
    wire N__44333;
    wire N__44332;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44318;
    wire N__44315;
    wire N__44314;
    wire N__44309;
    wire N__44308;
    wire N__44305;
    wire N__44302;
    wire N__44299;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44284;
    wire N__44281;
    wire N__44278;
    wire N__44273;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44252;
    wire N__44249;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44237;
    wire N__44234;
    wire N__44231;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44198;
    wire N__44195;
    wire N__44194;
    wire N__44193;
    wire N__44192;
    wire N__44189;
    wire N__44186;
    wire N__44183;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44171;
    wire N__44168;
    wire N__44165;
    wire N__44158;
    wire N__44153;
    wire N__44150;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44119;
    wire N__44116;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44101;
    wire N__44096;
    wire N__44093;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44082;
    wire N__44077;
    wire N__44074;
    wire N__44071;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44057;
    wire N__44056;
    wire N__44053;
    wire N__44050;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44036;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44024;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44014;
    wire N__44011;
    wire N__44008;
    wire N__44003;
    wire N__44000;
    wire N__43999;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43982;
    wire N__43979;
    wire N__43976;
    wire N__43975;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43958;
    wire N__43955;
    wire N__43952;
    wire N__43949;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43892;
    wire N__43889;
    wire N__43886;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43868;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43858;
    wire N__43855;
    wire N__43852;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43826;
    wire N__43823;
    wire N__43820;
    wire N__43817;
    wire N__43816;
    wire N__43813;
    wire N__43810;
    wire N__43805;
    wire N__43802;
    wire N__43799;
    wire N__43796;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43736;
    wire N__43733;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43676;
    wire N__43673;
    wire N__43670;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43637;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43627;
    wire N__43624;
    wire N__43621;
    wire N__43616;
    wire N__43613;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43586;
    wire N__43583;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43564;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43537;
    wire N__43534;
    wire N__43529;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43495;
    wire N__43492;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43475;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43463;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43412;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43397;
    wire N__43394;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43367;
    wire N__43364;
    wire N__43361;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43346;
    wire N__43343;
    wire N__43340;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43310;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43295;
    wire N__43292;
    wire N__43289;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43256;
    wire N__43253;
    wire N__43250;
    wire N__43247;
    wire N__43244;
    wire N__43241;
    wire N__43238;
    wire N__43235;
    wire N__43232;
    wire N__43229;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43214;
    wire N__43211;
    wire N__43208;
    wire N__43205;
    wire N__43202;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43184;
    wire N__43181;
    wire N__43178;
    wire N__43175;
    wire N__43172;
    wire N__43169;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43148;
    wire N__43145;
    wire N__43142;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43127;
    wire N__43124;
    wire N__43121;
    wire N__43118;
    wire N__43115;
    wire N__43112;
    wire N__43109;
    wire N__43108;
    wire N__43107;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43089;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43067;
    wire N__43066;
    wire N__43063;
    wire N__43060;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43022;
    wire N__43019;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42991;
    wire N__42988;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42975;
    wire N__42972;
    wire N__42969;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42947;
    wire N__42944;
    wire N__42943;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42927;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42880;
    wire N__42877;
    wire N__42876;
    wire N__42873;
    wire N__42870;
    wire N__42867;
    wire N__42864;
    wire N__42861;
    wire N__42858;
    wire N__42851;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42829;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42796;
    wire N__42793;
    wire N__42790;
    wire N__42787;
    wire N__42784;
    wire N__42779;
    wire N__42778;
    wire N__42777;
    wire N__42776;
    wire N__42775;
    wire N__42774;
    wire N__42773;
    wire N__42772;
    wire N__42771;
    wire N__42770;
    wire N__42769;
    wire N__42768;
    wire N__42767;
    wire N__42766;
    wire N__42765;
    wire N__42764;
    wire N__42763;
    wire N__42762;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42737;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42719;
    wire N__42716;
    wire N__42713;
    wire N__42712;
    wire N__42711;
    wire N__42710;
    wire N__42709;
    wire N__42708;
    wire N__42707;
    wire N__42706;
    wire N__42705;
    wire N__42704;
    wire N__42703;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42685;
    wire N__42676;
    wire N__42667;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42633;
    wire N__42632;
    wire N__42631;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42623;
    wire N__42622;
    wire N__42621;
    wire N__42620;
    wire N__42619;
    wire N__42618;
    wire N__42617;
    wire N__42616;
    wire N__42615;
    wire N__42614;
    wire N__42613;
    wire N__42608;
    wire N__42607;
    wire N__42606;
    wire N__42605;
    wire N__42602;
    wire N__42601;
    wire N__42600;
    wire N__42599;
    wire N__42598;
    wire N__42597;
    wire N__42596;
    wire N__42595;
    wire N__42586;
    wire N__42577;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42559;
    wire N__42556;
    wire N__42553;
    wire N__42552;
    wire N__42551;
    wire N__42550;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42542;
    wire N__42539;
    wire N__42538;
    wire N__42535;
    wire N__42534;
    wire N__42531;
    wire N__42530;
    wire N__42527;
    wire N__42526;
    wire N__42523;
    wire N__42522;
    wire N__42519;
    wire N__42518;
    wire N__42515;
    wire N__42514;
    wire N__42513;
    wire N__42510;
    wire N__42509;
    wire N__42506;
    wire N__42505;
    wire N__42502;
    wire N__42501;
    wire N__42498;
    wire N__42493;
    wire N__42490;
    wire N__42489;
    wire N__42488;
    wire N__42487;
    wire N__42486;
    wire N__42485;
    wire N__42484;
    wire N__42483;
    wire N__42482;
    wire N__42481;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42455;
    wire N__42454;
    wire N__42453;
    wire N__42452;
    wire N__42445;
    wire N__42440;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42428;
    wire N__42425;
    wire N__42424;
    wire N__42421;
    wire N__42420;
    wire N__42417;
    wire N__42416;
    wire N__42413;
    wire N__42396;
    wire N__42379;
    wire N__42364;
    wire N__42363;
    wire N__42362;
    wire N__42361;
    wire N__42360;
    wire N__42359;
    wire N__42358;
    wire N__42357;
    wire N__42356;
    wire N__42353;
    wire N__42348;
    wire N__42347;
    wire N__42346;
    wire N__42345;
    wire N__42344;
    wire N__42343;
    wire N__42342;
    wire N__42339;
    wire N__42330;
    wire N__42319;
    wire N__42316;
    wire N__42309;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42260;
    wire N__42251;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42226;
    wire N__42225;
    wire N__42224;
    wire N__42223;
    wire N__42222;
    wire N__42221;
    wire N__42220;
    wire N__42219;
    wire N__42218;
    wire N__42213;
    wire N__42212;
    wire N__42211;
    wire N__42206;
    wire N__42203;
    wire N__42202;
    wire N__42199;
    wire N__42198;
    wire N__42195;
    wire N__42194;
    wire N__42191;
    wire N__42190;
    wire N__42189;
    wire N__42182;
    wire N__42179;
    wire N__42174;
    wire N__42165;
    wire N__42162;
    wire N__42153;
    wire N__42144;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42110;
    wire N__42107;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42099;
    wire N__42098;
    wire N__42097;
    wire N__42096;
    wire N__42095;
    wire N__42092;
    wire N__42091;
    wire N__42086;
    wire N__42071;
    wire N__42068;
    wire N__42065;
    wire N__42062;
    wire N__42057;
    wire N__42048;
    wire N__42039;
    wire N__42034;
    wire N__42029;
    wire N__42026;
    wire N__42023;
    wire N__42020;
    wire N__42019;
    wire N__42016;
    wire N__42013;
    wire N__42008;
    wire N__42005;
    wire N__42004;
    wire N__42003;
    wire N__42002;
    wire N__42001;
    wire N__42000;
    wire N__41999;
    wire N__41998;
    wire N__41997;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41977;
    wire N__41974;
    wire N__41971;
    wire N__41966;
    wire N__41957;
    wire N__41950;
    wire N__41947;
    wire N__41944;
    wire N__41941;
    wire N__41936;
    wire N__41927;
    wire N__41916;
    wire N__41909;
    wire N__41906;
    wire N__41903;
    wire N__41896;
    wire N__41893;
    wire N__41888;
    wire N__41883;
    wire N__41880;
    wire N__41875;
    wire N__41870;
    wire N__41867;
    wire N__41864;
    wire N__41861;
    wire N__41858;
    wire N__41851;
    wire N__41842;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41821;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41801;
    wire N__41798;
    wire N__41795;
    wire N__41792;
    wire N__41789;
    wire N__41780;
    wire N__41777;
    wire N__41776;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41753;
    wire N__41750;
    wire N__41749;
    wire N__41746;
    wire N__41745;
    wire N__41742;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41728;
    wire N__41723;
    wire N__41722;
    wire N__41719;
    wire N__41718;
    wire N__41715;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41696;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41678;
    wire N__41675;
    wire N__41674;
    wire N__41671;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41657;
    wire N__41654;
    wire N__41649;
    wire N__41646;
    wire N__41639;
    wire N__41638;
    wire N__41635;
    wire N__41634;
    wire N__41631;
    wire N__41628;
    wire N__41625;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41600;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41561;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41540;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41528;
    wire N__41525;
    wire N__41522;
    wire N__41519;
    wire N__41516;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41504;
    wire N__41501;
    wire N__41498;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41486;
    wire N__41483;
    wire N__41480;
    wire N__41477;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41456;
    wire N__41453;
    wire N__41450;
    wire N__41447;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41429;
    wire N__41426;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41414;
    wire N__41411;
    wire N__41408;
    wire N__41405;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41300;
    wire N__41297;
    wire N__41294;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41273;
    wire N__41272;
    wire N__41269;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41255;
    wire N__41252;
    wire N__41247;
    wire N__41244;
    wire N__41237;
    wire N__41234;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41222;
    wire N__41219;
    wire N__41216;
    wire N__41213;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41165;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41140;
    wire N__41137;
    wire N__41134;
    wire N__41133;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41105;
    wire N__41104;
    wire N__41103;
    wire N__41100;
    wire N__41095;
    wire N__41094;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41078;
    wire N__41075;
    wire N__41074;
    wire N__41073;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41054;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41044;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41021;
    wire N__41020;
    wire N__41017;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40993;
    wire N__40990;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40957;
    wire N__40956;
    wire N__40955;
    wire N__40954;
    wire N__40951;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40941;
    wire N__40938;
    wire N__40937;
    wire N__40934;
    wire N__40931;
    wire N__40928;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40915;
    wire N__40912;
    wire N__40907;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40888;
    wire N__40885;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40862;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40851;
    wire N__40846;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40829;
    wire N__40826;
    wire N__40823;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40805;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40783;
    wire N__40780;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40763;
    wire N__40760;
    wire N__40757;
    wire N__40754;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40742;
    wire N__40739;
    wire N__40736;
    wire N__40735;
    wire N__40734;
    wire N__40729;
    wire N__40726;
    wire N__40721;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40709;
    wire N__40706;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40691;
    wire N__40688;
    wire N__40685;
    wire N__40682;
    wire N__40679;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40631;
    wire N__40630;
    wire N__40629;
    wire N__40628;
    wire N__40627;
    wire N__40626;
    wire N__40625;
    wire N__40624;
    wire N__40623;
    wire N__40622;
    wire N__40621;
    wire N__40620;
    wire N__40619;
    wire N__40618;
    wire N__40617;
    wire N__40616;
    wire N__40611;
    wire N__40610;
    wire N__40609;
    wire N__40608;
    wire N__40607;
    wire N__40606;
    wire N__40605;
    wire N__40604;
    wire N__40599;
    wire N__40594;
    wire N__40589;
    wire N__40584;
    wire N__40583;
    wire N__40582;
    wire N__40581;
    wire N__40580;
    wire N__40579;
    wire N__40578;
    wire N__40577;
    wire N__40568;
    wire N__40563;
    wire N__40560;
    wire N__40549;
    wire N__40544;
    wire N__40535;
    wire N__40526;
    wire N__40519;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40475;
    wire N__40474;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40454;
    wire N__40451;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40391;
    wire N__40388;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40370;
    wire N__40367;
    wire N__40364;
    wire N__40361;
    wire N__40358;
    wire N__40355;
    wire N__40352;
    wire N__40351;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40327;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40304;
    wire N__40301;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40286;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40273;
    wire N__40270;
    wire N__40267;
    wire N__40264;
    wire N__40259;
    wire N__40256;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40235;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40225;
    wire N__40222;
    wire N__40219;
    wire N__40216;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40136;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40103;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40085;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40070;
    wire N__40067;
    wire N__40064;
    wire N__40061;
    wire N__40058;
    wire N__40055;
    wire N__40052;
    wire N__40049;
    wire N__40046;
    wire N__40043;
    wire N__40040;
    wire N__40037;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40025;
    wire N__40022;
    wire N__40019;
    wire N__40016;
    wire N__40013;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__39998;
    wire N__39995;
    wire N__39992;
    wire N__39989;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39965;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39953;
    wire N__39950;
    wire N__39947;
    wire N__39944;
    wire N__39941;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39923;
    wire N__39920;
    wire N__39917;
    wire N__39914;
    wire N__39911;
    wire N__39908;
    wire N__39905;
    wire N__39902;
    wire N__39901;
    wire N__39898;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39877;
    wire N__39872;
    wire N__39871;
    wire N__39868;
    wire N__39865;
    wire N__39862;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39815;
    wire N__39812;
    wire N__39809;
    wire N__39806;
    wire N__39803;
    wire N__39800;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39778;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39755;
    wire N__39754;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39739;
    wire N__39738;
    wire N__39733;
    wire N__39730;
    wire N__39725;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39708;
    wire N__39703;
    wire N__39700;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39683;
    wire N__39682;
    wire N__39681;
    wire N__39678;
    wire N__39675;
    wire N__39672;
    wire N__39665;
    wire N__39664;
    wire N__39661;
    wire N__39660;
    wire N__39659;
    wire N__39658;
    wire N__39657;
    wire N__39656;
    wire N__39655;
    wire N__39654;
    wire N__39653;
    wire N__39652;
    wire N__39651;
    wire N__39650;
    wire N__39649;
    wire N__39648;
    wire N__39643;
    wire N__39640;
    wire N__39639;
    wire N__39638;
    wire N__39637;
    wire N__39636;
    wire N__39635;
    wire N__39634;
    wire N__39633;
    wire N__39628;
    wire N__39615;
    wire N__39606;
    wire N__39601;
    wire N__39586;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39578;
    wire N__39577;
    wire N__39574;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39555;
    wire N__39552;
    wire N__39539;
    wire N__39538;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39528;
    wire N__39525;
    wire N__39522;
    wire N__39515;
    wire N__39514;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39496;
    wire N__39495;
    wire N__39490;
    wire N__39487;
    wire N__39482;
    wire N__39481;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39463;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39451;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39436;
    wire N__39431;
    wire N__39430;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39419;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39405;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39389;
    wire N__39386;
    wire N__39385;
    wire N__39382;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39364;
    wire N__39363;
    wire N__39358;
    wire N__39355;
    wire N__39350;
    wire N__39349;
    wire N__39348;
    wire N__39343;
    wire N__39340;
    wire N__39339;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39322;
    wire N__39317;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39301;
    wire N__39298;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39281;
    wire N__39280;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39254;
    wire N__39251;
    wire N__39242;
    wire N__39241;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39223;
    wire N__39218;
    wire N__39215;
    wire N__39214;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39191;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39179;
    wire N__39178;
    wire N__39175;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39149;
    wire N__39148;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39130;
    wire N__39129;
    wire N__39124;
    wire N__39121;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39107;
    wire N__39104;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39087;
    wire N__39080;
    wire N__39079;
    wire N__39078;
    wire N__39077;
    wire N__39076;
    wire N__39075;
    wire N__39074;
    wire N__39059;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39011;
    wire N__39010;
    wire N__39007;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38990;
    wire N__38989;
    wire N__38988;
    wire N__38983;
    wire N__38980;
    wire N__38975;
    wire N__38974;
    wire N__38971;
    wire N__38966;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38936;
    wire N__38935;
    wire N__38930;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38906;
    wire N__38903;
    wire N__38902;
    wire N__38901;
    wire N__38896;
    wire N__38893;
    wire N__38888;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38870;
    wire N__38867;
    wire N__38866;
    wire N__38865;
    wire N__38860;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38821;
    wire N__38818;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38794;
    wire N__38791;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38752;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38683;
    wire N__38680;
    wire N__38677;
    wire N__38674;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38659;
    wire N__38656;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38629;
    wire N__38626;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38608;
    wire N__38605;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38570;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38558;
    wire N__38555;
    wire N__38552;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38534;
    wire N__38533;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38513;
    wire N__38512;
    wire N__38509;
    wire N__38506;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38426;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38411;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38399;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38387;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38375;
    wire N__38372;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38342;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38334;
    wire N__38331;
    wire N__38326;
    wire N__38323;
    wire N__38318;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38293;
    wire N__38288;
    wire N__38287;
    wire N__38282;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38262;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38248;
    wire N__38243;
    wire N__38242;
    wire N__38239;
    wire N__38238;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38219;
    wire N__38216;
    wire N__38215;
    wire N__38214;
    wire N__38211;
    wire N__38208;
    wire N__38205;
    wire N__38200;
    wire N__38195;
    wire N__38194;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38182;
    wire N__38179;
    wire N__38174;
    wire N__38173;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38147;
    wire N__38146;
    wire N__38141;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38129;
    wire N__38126;
    wire N__38125;
    wire N__38124;
    wire N__38121;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38096;
    wire N__38093;
    wire N__38092;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38075;
    wire N__38072;
    wire N__38069;
    wire N__38066;
    wire N__38063;
    wire N__38060;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38038;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38023;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38006;
    wire N__38003;
    wire N__38000;
    wire N__37999;
    wire N__37996;
    wire N__37995;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37979;
    wire N__37976;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37955;
    wire N__37952;
    wire N__37949;
    wire N__37946;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37874;
    wire N__37871;
    wire N__37868;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37822;
    wire N__37821;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37805;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37778;
    wire N__37775;
    wire N__37772;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37735;
    wire N__37732;
    wire N__37731;
    wire N__37730;
    wire N__37729;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37698;
    wire N__37685;
    wire N__37682;
    wire N__37681;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37658;
    wire N__37655;
    wire N__37652;
    wire N__37649;
    wire N__37648;
    wire N__37647;
    wire N__37644;
    wire N__37643;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37635;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37600;
    wire N__37595;
    wire N__37590;
    wire N__37587;
    wire N__37582;
    wire N__37579;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37484;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37472;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37438;
    wire N__37435;
    wire N__37432;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37293;
    wire N__37288;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37277;
    wire N__37276;
    wire N__37273;
    wire N__37270;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37250;
    wire N__37249;
    wire N__37244;
    wire N__37243;
    wire N__37242;
    wire N__37239;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37211;
    wire N__37206;
    wire N__37199;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36920;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36898;
    wire N__36897;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36886;
    wire N__36885;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36871;
    wire N__36870;
    wire N__36867;
    wire N__36866;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36845;
    wire N__36842;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36812;
    wire N__36809;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36589;
    wire N__36584;
    wire N__36583;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36556;
    wire N__36553;
    wire N__36550;
    wire N__36545;
    wire N__36542;
    wire N__36541;
    wire N__36538;
    wire N__36535;
    wire N__36530;
    wire N__36527;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36515;
    wire N__36512;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36460;
    wire N__36457;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36434;
    wire N__36431;
    wire N__36430;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36414;
    wire N__36407;
    wire N__36406;
    wire N__36405;
    wire N__36398;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36356;
    wire N__36353;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36341;
    wire N__36338;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36326;
    wire N__36323;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36302;
    wire N__36299;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36287;
    wire N__36284;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36272;
    wire N__36269;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36257;
    wire N__36254;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36242;
    wire N__36239;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36227;
    wire N__36224;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36212;
    wire N__36209;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36197;
    wire N__36194;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36182;
    wire N__36179;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36143;
    wire N__36140;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36128;
    wire N__36125;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36113;
    wire N__36110;
    wire N__36109;
    wire N__36106;
    wire N__36103;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36064;
    wire N__36061;
    wire N__36058;
    wire N__36053;
    wire N__36050;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36038;
    wire N__36035;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36023;
    wire N__36020;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36008;
    wire N__36005;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35986;
    wire N__35985;
    wire N__35984;
    wire N__35983;
    wire N__35982;
    wire N__35981;
    wire N__35980;
    wire N__35977;
    wire N__35974;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35963;
    wire N__35962;
    wire N__35959;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35947;
    wire N__35936;
    wire N__35927;
    wire N__35924;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35876;
    wire N__35873;
    wire N__35870;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35819;
    wire N__35816;
    wire N__35813;
    wire N__35810;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35663;
    wire N__35662;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35645;
    wire N__35642;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35632;
    wire N__35627;
    wire N__35624;
    wire N__35623;
    wire N__35622;
    wire N__35621;
    wire N__35620;
    wire N__35619;
    wire N__35618;
    wire N__35617;
    wire N__35616;
    wire N__35615;
    wire N__35614;
    wire N__35613;
    wire N__35612;
    wire N__35611;
    wire N__35610;
    wire N__35609;
    wire N__35608;
    wire N__35607;
    wire N__35606;
    wire N__35605;
    wire N__35604;
    wire N__35603;
    wire N__35602;
    wire N__35601;
    wire N__35600;
    wire N__35599;
    wire N__35590;
    wire N__35589;
    wire N__35588;
    wire N__35587;
    wire N__35586;
    wire N__35581;
    wire N__35572;
    wire N__35563;
    wire N__35554;
    wire N__35545;
    wire N__35536;
    wire N__35533;
    wire N__35524;
    wire N__35519;
    wire N__35510;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35483;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35459;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35441;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35257;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35247;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35233;
    wire N__35232;
    wire N__35229;
    wire N__35226;
    wire N__35223;
    wire N__35216;
    wire N__35213;
    wire N__35210;
    wire N__35209;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35199;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35185;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35161;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35137;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35113;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35096;
    wire N__35093;
    wire N__35092;
    wire N__35091;
    wire N__35088;
    wire N__35083;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35071;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35047;
    wire N__35046;
    wire N__35043;
    wire N__35040;
    wire N__35037;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35023;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35013;
    wire N__35006;
    wire N__35003;
    wire N__35000;
    wire N__34999;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34975;
    wire N__34974;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34951;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34927;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34903;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34886;
    wire N__34883;
    wire N__34882;
    wire N__34881;
    wire N__34878;
    wire N__34873;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34861;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34844;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34825;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34813;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34789;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34765;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34741;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34717;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34700;
    wire N__34697;
    wire N__34694;
    wire N__34693;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34658;
    wire N__34657;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34625;
    wire N__34624;
    wire N__34619;
    wire N__34616;
    wire N__34615;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34592;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34577;
    wire N__34576;
    wire N__34571;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34556;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34546;
    wire N__34545;
    wire N__34544;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34527;
    wire N__34524;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34506;
    wire N__34503;
    wire N__34496;
    wire N__34495;
    wire N__34494;
    wire N__34493;
    wire N__34492;
    wire N__34491;
    wire N__34490;
    wire N__34489;
    wire N__34488;
    wire N__34487;
    wire N__34486;
    wire N__34485;
    wire N__34484;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34472;
    wire N__34463;
    wire N__34462;
    wire N__34461;
    wire N__34460;
    wire N__34459;
    wire N__34458;
    wire N__34457;
    wire N__34456;
    wire N__34455;
    wire N__34446;
    wire N__34437;
    wire N__34436;
    wire N__34435;
    wire N__34434;
    wire N__34433;
    wire N__34428;
    wire N__34421;
    wire N__34410;
    wire N__34409;
    wire N__34408;
    wire N__34407;
    wire N__34406;
    wire N__34401;
    wire N__34392;
    wire N__34387;
    wire N__34384;
    wire N__34375;
    wire N__34366;
    wire N__34361;
    wire N__34360;
    wire N__34359;
    wire N__34358;
    wire N__34355;
    wire N__34348;
    wire N__34345;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34310;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34274;
    wire N__34271;
    wire N__34270;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34260;
    wire N__34259;
    wire N__34256;
    wire N__34251;
    wire N__34248;
    wire N__34247;
    wire N__34246;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34198;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34181;
    wire N__34178;
    wire N__34175;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34167;
    wire N__34162;
    wire N__34159;
    wire N__34154;
    wire N__34153;
    wire N__34150;
    wire N__34145;
    wire N__34144;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34129;
    wire N__34124;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34102;
    wire N__34097;
    wire N__34094;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34086;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34063;
    wire N__34062;
    wire N__34061;
    wire N__34058;
    wire N__34051;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34023;
    wire N__34022;
    wire N__34021;
    wire N__34018;
    wire N__34017;
    wire N__34014;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33965;
    wire N__33964;
    wire N__33959;
    wire N__33956;
    wire N__33955;
    wire N__33950;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33935;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33923;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33833;
    wire N__33830;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33755;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33743;
    wire N__33742;
    wire N__33737;
    wire N__33734;
    wire N__33733;
    wire N__33730;
    wire N__33727;
    wire N__33722;
    wire N__33719;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33707;
    wire N__33704;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33671;
    wire N__33668;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33521;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33376;
    wire N__33375;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33356;
    wire N__33353;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33226;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33050;
    wire N__33047;
    wire N__33046;
    wire N__33041;
    wire N__33038;
    wire N__33035;
    wire N__33032;
    wire N__33029;
    wire N__33026;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32939;
    wire N__32936;
    wire N__32933;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32840;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32725;
    wire N__32722;
    wire N__32719;
    wire N__32716;
    wire N__32713;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32698;
    wire N__32695;
    wire N__32692;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32677;
    wire N__32676;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32655;
    wire N__32652;
    wire N__32647;
    wire N__32644;
    wire N__32639;
    wire N__32638;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32608;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32588;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32527;
    wire N__32524;
    wire N__32519;
    wire N__32516;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32486;
    wire N__32483;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32471;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32456;
    wire N__32453;
    wire N__32452;
    wire N__32447;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32432;
    wire N__32429;
    wire N__32428;
    wire N__32425;
    wire N__32422;
    wire N__32417;
    wire N__32416;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32402;
    wire N__32399;
    wire N__32398;
    wire N__32393;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32383;
    wire N__32378;
    wire N__32375;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32367;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32351;
    wire N__32348;
    wire N__32347;
    wire N__32346;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32330;
    wire N__32327;
    wire N__32326;
    wire N__32321;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32306;
    wire N__32303;
    wire N__32302;
    wire N__32297;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32287;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32261;
    wire N__32258;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32243;
    wire N__32240;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32213;
    wire N__32210;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32198;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32183;
    wire N__32180;
    wire N__32179;
    wire N__32174;
    wire N__32171;
    wire N__32170;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32156;
    wire N__32153;
    wire N__32152;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32117;
    wire N__32114;
    wire N__32113;
    wire N__32110;
    wire N__32107;
    wire N__32104;
    wire N__32099;
    wire N__32096;
    wire N__32095;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32081;
    wire N__32078;
    wire N__32077;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32042;
    wire N__32039;
    wire N__32038;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32017;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31969;
    wire N__31964;
    wire N__31961;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31946;
    wire N__31943;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31907;
    wire N__31904;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31786;
    wire N__31785;
    wire N__31782;
    wire N__31781;
    wire N__31780;
    wire N__31779;
    wire N__31778;
    wire N__31775;
    wire N__31774;
    wire N__31773;
    wire N__31772;
    wire N__31771;
    wire N__31770;
    wire N__31769;
    wire N__31768;
    wire N__31767;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31759;
    wire N__31758;
    wire N__31757;
    wire N__31756;
    wire N__31747;
    wire N__31744;
    wire N__31737;
    wire N__31736;
    wire N__31735;
    wire N__31734;
    wire N__31733;
    wire N__31732;
    wire N__31731;
    wire N__31730;
    wire N__31729;
    wire N__31728;
    wire N__31727;
    wire N__31720;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31698;
    wire N__31693;
    wire N__31690;
    wire N__31685;
    wire N__31682;
    wire N__31677;
    wire N__31668;
    wire N__31665;
    wire N__31660;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31490;
    wire N__31487;
    wire N__31484;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31381;
    wire N__31376;
    wire N__31373;
    wire N__31372;
    wire N__31367;
    wire N__31364;
    wire N__31363;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31315;
    wire N__31310;
    wire N__31307;
    wire N__31306;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31294;
    wire N__31289;
    wire N__31286;
    wire N__31285;
    wire N__31280;
    wire N__31277;
    wire N__31276;
    wire N__31271;
    wire N__31268;
    wire N__31267;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31255;
    wire N__31250;
    wire N__31247;
    wire N__31246;
    wire N__31241;
    wire N__31238;
    wire N__31235;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31220;
    wire N__31219;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31123;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31097;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30874;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30811;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30730;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30722;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30685;
    wire N__30684;
    wire N__30683;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30675;
    wire N__30672;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30638;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30623;
    wire N__30620;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30584;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30488;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30466;
    wire N__30461;
    wire N__30458;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30443;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30432;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30367;
    wire N__30364;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30347;
    wire N__30344;
    wire N__30343;
    wire N__30340;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30317;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30224;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30206;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29879;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29774;
    wire N__29773;
    wire N__29772;
    wire N__29771;
    wire N__29764;
    wire N__29761;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29716;
    wire N__29715;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29699;
    wire N__29698;
    wire N__29693;
    wire N__29690;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29682;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29666;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29651;
    wire N__29650;
    wire N__29649;
    wire N__29648;
    wire N__29639;
    wire N__29636;
    wire N__29633;
    wire N__29630;
    wire N__29629;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29614;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29597;
    wire N__29594;
    wire N__29593;
    wire N__29592;
    wire N__29587;
    wire N__29584;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29566;
    wire N__29565;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29549;
    wire N__29548;
    wire N__29547;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29531;
    wire N__29530;
    wire N__29529;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29513;
    wire N__29512;
    wire N__29511;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29495;
    wire N__29492;
    wire N__29491;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29476;
    wire N__29471;
    wire N__29468;
    wire N__29467;
    wire N__29464;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29441;
    wire N__29440;
    wire N__29439;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29423;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29415;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29392;
    wire N__29391;
    wire N__29390;
    wire N__29389;
    wire N__29388;
    wire N__29387;
    wire N__29386;
    wire N__29385;
    wire N__29384;
    wire N__29383;
    wire N__29382;
    wire N__29381;
    wire N__29380;
    wire N__29379;
    wire N__29378;
    wire N__29369;
    wire N__29360;
    wire N__29359;
    wire N__29358;
    wire N__29357;
    wire N__29356;
    wire N__29355;
    wire N__29354;
    wire N__29353;
    wire N__29352;
    wire N__29351;
    wire N__29350;
    wire N__29349;
    wire N__29348;
    wire N__29347;
    wire N__29346;
    wire N__29345;
    wire N__29344;
    wire N__29337;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29311;
    wire N__29302;
    wire N__29293;
    wire N__29284;
    wire N__29279;
    wire N__29264;
    wire N__29261;
    wire N__29260;
    wire N__29257;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29249;
    wire N__29246;
    wire N__29241;
    wire N__29238;
    wire N__29233;
    wire N__29230;
    wire N__29225;
    wire N__29224;
    wire N__29223;
    wire N__29220;
    wire N__29215;
    wire N__29210;
    wire N__29209;
    wire N__29208;
    wire N__29205;
    wire N__29200;
    wire N__29195;
    wire N__29194;
    wire N__29193;
    wire N__29190;
    wire N__29185;
    wire N__29180;
    wire N__29179;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29162;
    wire N__29161;
    wire N__29160;
    wire N__29155;
    wire N__29152;
    wire N__29149;
    wire N__29144;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29136;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29019;
    wire N__29016;
    wire N__29011;
    wire N__29008;
    wire N__29003;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28987;
    wire N__28986;
    wire N__28983;
    wire N__28978;
    wire N__28973;
    wire N__28972;
    wire N__28969;
    wire N__28968;
    wire N__28967;
    wire N__28962;
    wire N__28957;
    wire N__28954;
    wire N__28949;
    wire N__28946;
    wire N__28943;
    wire N__28942;
    wire N__28941;
    wire N__28938;
    wire N__28933;
    wire N__28928;
    wire N__28925;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28912;
    wire N__28909;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28892;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28880;
    wire N__28879;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28867;
    wire N__28862;
    wire N__28861;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28837;
    wire N__28836;
    wire N__28835;
    wire N__28834;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28830;
    wire N__28829;
    wire N__28828;
    wire N__28827;
    wire N__28818;
    wire N__28817;
    wire N__28816;
    wire N__28815;
    wire N__28814;
    wire N__28813;
    wire N__28812;
    wire N__28811;
    wire N__28810;
    wire N__28809;
    wire N__28808;
    wire N__28807;
    wire N__28806;
    wire N__28797;
    wire N__28788;
    wire N__28787;
    wire N__28786;
    wire N__28785;
    wire N__28784;
    wire N__28783;
    wire N__28782;
    wire N__28781;
    wire N__28780;
    wire N__28777;
    wire N__28768;
    wire N__28759;
    wire N__28750;
    wire N__28745;
    wire N__28736;
    wire N__28727;
    wire N__28722;
    wire N__28715;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28699;
    wire N__28696;
    wire N__28695;
    wire N__28692;
    wire N__28691;
    wire N__28688;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28640;
    wire N__28639;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28619;
    wire N__28618;
    wire N__28615;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28567;
    wire N__28562;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28547;
    wire N__28546;
    wire N__28545;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28499;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28451;
    wire N__28450;
    wire N__28449;
    wire N__28446;
    wire N__28441;
    wire N__28436;
    wire N__28435;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28412;
    wire N__28409;
    wire N__28408;
    wire N__28407;
    wire N__28404;
    wire N__28399;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28369;
    wire N__28364;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28352;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27830;
    wire N__27827;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27722;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27682;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27632;
    wire N__27629;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27578;
    wire N__27575;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27494;
    wire N__27491;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27479;
    wire N__27476;
    wire N__27475;
    wire N__27472;
    wire N__27469;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27434;
    wire N__27431;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27323;
    wire N__27320;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27287;
    wire N__27284;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27272;
    wire N__27269;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27224;
    wire N__27221;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27149;
    wire N__27146;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27113;
    wire N__27110;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27098;
    wire N__27095;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27073;
    wire N__27068;
    wire N__27065;
    wire N__27064;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26981;
    wire N__26980;
    wire N__26977;
    wire N__26976;
    wire N__26975;
    wire N__26972;
    wire N__26971;
    wire N__26970;
    wire N__26969;
    wire N__26966;
    wire N__26961;
    wire N__26958;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26910;
    wire N__26907;
    wire N__26902;
    wire N__26899;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26884;
    wire N__26883;
    wire N__26880;
    wire N__26875;
    wire N__26870;
    wire N__26867;
    wire N__26866;
    wire N__26865;
    wire N__26862;
    wire N__26855;
    wire N__26852;
    wire N__26851;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26803;
    wire N__26798;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26787;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26759;
    wire N__26758;
    wire N__26753;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26731;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26723;
    wire N__26716;
    wire N__26713;
    wire N__26708;
    wire N__26707;
    wire N__26706;
    wire N__26705;
    wire N__26704;
    wire N__26699;
    wire N__26698;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26678;
    wire N__26677;
    wire N__26676;
    wire N__26673;
    wire N__26668;
    wire N__26665;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26653;
    wire N__26652;
    wire N__26651;
    wire N__26644;
    wire N__26641;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26626;
    wire N__26625;
    wire N__26624;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26599;
    wire N__26596;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26576;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26502;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26486;
    wire N__26483;
    wire N__26482;
    wire N__26481;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26312;
    wire N__26309;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26207;
    wire N__26204;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26189;
    wire N__26186;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26156;
    wire N__26153;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26030;
    wire N__26027;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25930;
    wire N__25925;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25910;
    wire N__25907;
    wire N__25906;
    wire N__25901;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25876;
    wire N__25875;
    wire N__25874;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25866;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25829;
    wire N__25828;
    wire N__25823;
    wire N__25820;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25808;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25447;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25433;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25348;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25285;
    wire N__25284;
    wire N__25283;
    wire N__25282;
    wire N__25281;
    wire N__25280;
    wire N__25279;
    wire N__25278;
    wire N__25277;
    wire N__25276;
    wire N__25275;
    wire N__25274;
    wire N__25273;
    wire N__25272;
    wire N__25271;
    wire N__25270;
    wire N__25269;
    wire N__25268;
    wire N__25267;
    wire N__25266;
    wire N__25265;
    wire N__25264;
    wire N__25263;
    wire N__25262;
    wire N__25261;
    wire N__25260;
    wire N__25259;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25255;
    wire N__25246;
    wire N__25237;
    wire N__25228;
    wire N__25219;
    wire N__25210;
    wire N__25201;
    wire N__25192;
    wire N__25183;
    wire N__25176;
    wire N__25163;
    wire N__25160;
    wire N__25159;
    wire N__25158;
    wire N__25157;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24961;
    wire N__24960;
    wire N__24957;
    wire N__24952;
    wire N__24947;
    wire N__24944;
    wire N__24943;
    wire N__24942;
    wire N__24939;
    wire N__24934;
    wire N__24929;
    wire N__24926;
    wire N__24925;
    wire N__24924;
    wire N__24921;
    wire N__24916;
    wire N__24911;
    wire N__24908;
    wire N__24907;
    wire N__24906;
    wire N__24903;
    wire N__24898;
    wire N__24893;
    wire N__24890;
    wire N__24889;
    wire N__24888;
    wire N__24885;
    wire N__24880;
    wire N__24875;
    wire N__24872;
    wire N__24871;
    wire N__24870;
    wire N__24867;
    wire N__24862;
    wire N__24857;
    wire N__24854;
    wire N__24853;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24838;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24803;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24788;
    wire N__24785;
    wire N__24784;
    wire N__24779;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24764;
    wire N__24761;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24749;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24734;
    wire N__24731;
    wire N__24730;
    wire N__24725;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24710;
    wire N__24707;
    wire N__24706;
    wire N__24705;
    wire N__24702;
    wire N__24697;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24652;
    wire N__24651;
    wire N__24644;
    wire N__24641;
    wire N__24640;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24626;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24620;
    wire N__24619;
    wire N__24616;
    wire N__24615;
    wire N__24612;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24584;
    wire N__24583;
    wire N__24582;
    wire N__24577;
    wire N__24574;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24556;
    wire N__24551;
    wire N__24548;
    wire N__24547;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24523;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24511;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24496;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24457;
    wire N__24456;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24448;
    wire N__24447;
    wire N__24444;
    wire N__24443;
    wire N__24440;
    wire N__24439;
    wire N__24438;
    wire N__24437;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24407;
    wire N__24406;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24387;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24365;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24335;
    wire N__24334;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24322;
    wire N__24319;
    wire N__24316;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24304;
    wire N__24299;
    wire N__24296;
    wire N__24295;
    wire N__24290;
    wire N__24287;
    wire N__24286;
    wire N__24281;
    wire N__24278;
    wire N__24277;
    wire N__24272;
    wire N__24269;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24232;
    wire N__24227;
    wire N__24224;
    wire N__24223;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24184;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24164;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24127;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24091;
    wire N__24088;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24052;
    wire N__24049;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23902;
    wire N__23901;
    wire N__23900;
    wire N__23899;
    wire N__23890;
    wire N__23889;
    wire N__23886;
    wire N__23885;
    wire N__23884;
    wire N__23881;
    wire N__23880;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23868;
    wire N__23865;
    wire N__23860;
    wire N__23857;
    wire N__23852;
    wire N__23849;
    wire N__23844;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23785;
    wire N__23782;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23758;
    wire N__23755;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23707;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23677;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23632;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23590;
    wire N__23589;
    wire N__23588;
    wire N__23587;
    wire N__23586;
    wire N__23585;
    wire N__23584;
    wire N__23583;
    wire N__23582;
    wire N__23573;
    wire N__23568;
    wire N__23559;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23525;
    wire N__23522;
    wire N__23521;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23494;
    wire N__23493;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23485;
    wire N__23482;
    wire N__23481;
    wire N__23478;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23344;
    wire N__23341;
    wire N__23338;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23234;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23195;
    wire N__23194;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23149;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire \pwm_generator_inst.O_0_1 ;
    wire \pwm_generator_inst.O_0_0 ;
    wire \pwm_generator_inst.O_0_5 ;
    wire \pwm_generator_inst.O_0_3 ;
    wire \pwm_generator_inst.O_0_4 ;
    wire \pwm_generator_inst.O_0_2 ;
    wire \pwm_generator_inst.O_0_6 ;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_0 ;
    wire bfn_1_13_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_8 ;
    wire bfn_1_14_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_8 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_9 ;
    wire \pwm_generator_inst.O_11 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_11 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_10 ;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_11 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_12 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_15 ;
    wire bfn_1_15_0_;
    wire \pwm_generator_inst.un18_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_18 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_19 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_20 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_21 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_22 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_23 ;
    wire bfn_1_16_0_;
    wire \pwm_generator_inst.un18_threshold_1_cry_24 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_25 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_20 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_22 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_21 ;
    wire \pwm_generator_inst.un5_threshold_2_0 ;
    wire \pwm_generator_inst.un5_threshold_1_15 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_15 ;
    wire bfn_1_17_0_;
    wire \pwm_generator_inst.un5_threshold_2_1 ;
    wire \pwm_generator_inst.un5_threshold_1_16 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un5_threshold_2_2 ;
    wire \pwm_generator_inst.un5_threshold_1_17 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un5_threshold_2_3 ;
    wire \pwm_generator_inst.un5_threshold_1_18 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un5_threshold_2_4 ;
    wire \pwm_generator_inst.un5_threshold_1_19 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un5_threshold_2_5 ;
    wire \pwm_generator_inst.un5_threshold_1_20 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un5_threshold_1_21 ;
    wire \pwm_generator_inst.un5_threshold_2_6 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un5_threshold_1_22 ;
    wire \pwm_generator_inst.un5_threshold_2_7 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un5_threshold_1_23 ;
    wire \pwm_generator_inst.un5_threshold_2_8 ;
    wire bfn_1_18_0_;
    wire \pwm_generator_inst.un5_threshold_1_24 ;
    wire \pwm_generator_inst.un5_threshold_2_9 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un5_threshold_1_25 ;
    wire \pwm_generator_inst.un5_threshold_2_10 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un5_threshold_2_11 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un5_threshold_2_12 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un5_threshold_2_13 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un5_threshold_2_14 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_15 ;
    wire bfn_1_19_0_;
    wire bfn_1_20_0_;
    wire \pwm_generator_inst.O_0_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_0_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_0_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.O_0_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.O_0_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.O_0_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.O_0_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0 ;
    wire bfn_1_21_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8 ;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7 ;
    wire bfn_1_22_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0 ;
    wire N_112_i_i;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0 ;
    wire \pwm_generator_inst.un1_counterlto2_0 ;
    wire bfn_2_15_0_;
    wire \pwm_generator_inst.un18_threshold1_18 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1_cry_0 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_1 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_2 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_3 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_4 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_5 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_7 ;
    wire bfn_2_16_0_;
    wire \pwm_generator_inst.un22_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO ;
    wire \pwm_generator_inst.un18_threshold1_25 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO ;
    wire \pwm_generator_inst.un18_threshold1_23 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_23 ;
    wire \pwm_generator_inst.un18_threshold1_24 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_24 ;
    wire \pwm_generator_inst.un5_threshold_1_26 ;
    wire \pwm_generator_inst.un5_threshold_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_ ;
    wire \pwm_generator_inst.un5_threshold_2_1_15 ;
    wire \pwm_generator_inst.un5_threshold_add_1_axb_16 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_25 ;
    wire un8_start_stop;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire bfn_3_12_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_3_13_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO ;
    wire \pwm_generator_inst.un18_threshold1_19 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_19 ;
    wire \pwm_generator_inst.un18_threshold1_20 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO ;
    wire \pwm_generator_inst.un18_threshold1_21 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1 ;
    wire \pwm_generator_inst.un18_threshold1_22 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0 ;
    wire \pwm_generator_inst.N_179_i ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_3_15_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.N_180_i ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.N_181_i ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.N_182_i ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.N_183_i ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.N_184_i ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.N_185_i ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.N_186_i ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.N_187_i ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_3_16_0_;
    wire \pwm_generator_inst.N_188_i ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31_cascade_;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire elapsed_time_ns_1_RNI1BOBB_0_14_cascade_;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_start_0 ;
    wire \phase_controller_inst2.stateZ0Z_4 ;
    wire \phase_controller_inst2.start_flagZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire bfn_8_8_0_;
    wire \phase_controller_inst2.stoper_tr.counter_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_7 ;
    wire bfn_8_9_0_;
    wire \phase_controller_inst2.stoper_tr.counter_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_16 ;
    wire bfn_8_10_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_23 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_24 ;
    wire bfn_8_11_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_i_0 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0_g ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_0 ;
    wire bfn_8_12_0_;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_1 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_8 ;
    wire bfn_8_13_0_;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_9 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ;
    wire bfn_8_14_0_;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_30 ;
    wire bfn_8_15_0_;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.counter ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire elapsed_time_ns_1_RNI2COBB_0_15_cascade_;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ;
    wire bfn_8_16_0_;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_1;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_2;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_3;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_4;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_5;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_6;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_7;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_8;
    wire bfn_8_17_0_;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_9;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_10;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_11;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_12;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_13;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_14;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_15;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_16;
    wire bfn_8_18_0_;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_17;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_18;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_19;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ;
    wire bfn_8_19_0_;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_27;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ;
    wire bfn_8_20_0_;
    wire \phase_controller_inst1.stoper_tr.counter_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_7 ;
    wire bfn_8_21_0_;
    wire \phase_controller_inst1.stoper_tr.counter_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_15 ;
    wire bfn_8_22_0_;
    wire \phase_controller_inst1.stoper_tr.counter_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_23 ;
    wire bfn_8_23_0_;
    wire \phase_controller_inst1.stoper_tr.counter_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0_g ;
    wire s4_phy_c;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.state_ns_0_0_1 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire il_max_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.un4_start_0 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire start_stop_c;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.state_ns_0_0_1_cascade_ ;
    wire \phase_controller_inst1.start_flagZ0 ;
    wire \phase_controller_inst1.stoper_tr.un4_start_0_cascade_ ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire elapsed_time_ns_1_RNIJI91B_0_7_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire elapsed_time_ns_1_RNIFE91B_0_3_cascade_;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ;
    wire bfn_9_14_0_;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ;
    wire bfn_9_15_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ;
    wire bfn_9_16_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ;
    wire bfn_9_17_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_28;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_0 ;
    wire bfn_9_18_0_;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_1 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_8 ;
    wire bfn_9_19_0_;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_9 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ;
    wire bfn_9_20_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_30 ;
    wire bfn_9_21_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.counter ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_24;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_25;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt26 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_26;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_i_0 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire s3_phy_c;
    wire bfn_10_2_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_7 ;
    wire bfn_10_3_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_15 ;
    wire bfn_10_4_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_23 ;
    wire bfn_10_5_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_i_0 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ;
    wire il_min_comp1_c;
    wire il_max_comp1_c;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire elapsed_time_ns_1_RNI0AOBB_0_13_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire elapsed_time_ns_1_RNIKJ91B_0_8_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire \pwm_generator_inst.un3_threshold_iZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire elapsed_time_ns_1_RNIIH91B_0_6_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire elapsed_time_ns_1_RNILK91B_0_9_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire elapsed_time_ns_1_RNIGF91B_0_4_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire elapsed_time_ns_1_RNIU8PBB_0_20_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire elapsed_time_ns_1_RNIHG91B_0_5_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire elapsed_time_ns_1_RNI3DOBB_0_16_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire elapsed_time_ns_1_RNIT6OBB_0_10_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire elapsed_time_ns_1_RNI4EOBB_0_17_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire elapsed_time_ns_1_RNI4FPBB_0_26_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire elapsed_time_ns_1_RNI5FOBB_0_18_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire elapsed_time_ns_1_RNI5GPBB_0_27_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire elapsed_time_ns_1_RNI3EPBB_0_25_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire elapsed_time_ns_1_RNI6HPBB_0_28_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_20;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_21;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_22;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_23;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt20 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire elapsed_time_ns_1_RNI6GOBB_0_19_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.counter ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_0 ;
    wire bfn_11_4_0_;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_1 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_8 ;
    wire bfn_11_5_0_;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_9 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ;
    wire bfn_11_6_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt30 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_30 ;
    wire bfn_11_7_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_0 ;
    wire bfn_11_12_0_;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_8 ;
    wire bfn_11_13_0_;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_15 ;
    wire bfn_11_14_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_30 ;
    wire bfn_11_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire elapsed_time_ns_1_RNI0BPBB_0_22_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.counter ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_0 ;
    wire bfn_11_16_0_;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_8 ;
    wire bfn_11_17_0_;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_15 ;
    wire bfn_11_18_0_;
    wire \phase_controller_inst1.stoper_hc.counter_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_24 ;
    wire bfn_11_19_0_;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire bfn_11_20_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire bfn_11_21_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire bfn_11_22_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_11_23_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ;
    wire bfn_12_7_0_;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_1;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_5;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_8;
    wire bfn_12_8_0_;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_9;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_11;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_12;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_13;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_14;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_15;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ;
    wire bfn_12_9_0_;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_20;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_21;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_22;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_23;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_24;
    wire bfn_12_10_0_;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_26;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_27;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_4;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_2;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_6;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_19;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_3;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_7;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_10;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_25;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.N_167_i ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt16 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_16;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_17;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt18 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_18;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_i_0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_12_19_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_12_20_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_12_21_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_12_22_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_168_i ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_12_23_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_12_24_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire GB_BUFFER_red_c_g_THRU_CO;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire elapsed_time_ns_1_RNI24CN9_0_15_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ;
    wire bfn_13_7_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ;
    wire bfn_13_8_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ;
    wire bfn_13_9_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ;
    wire bfn_13_10_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_28;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt30 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_8 ;
    wire bfn_13_21_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ;
    wire bfn_13_22_0_;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire elapsed_time_ns_1_RNITUBN9_0_10_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire elapsed_time_ns_1_RNIUVBN9_0_11_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire elapsed_time_ns_1_RNIJ53T9_0_7_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire elapsed_time_ns_1_RNIK63T9_0_8_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire elapsed_time_ns_1_RNI47DN9_0_26_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire elapsed_time_ns_1_RNIL73T9_0_9_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire elapsed_time_ns_1_RNI14DN9_0_23_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire elapsed_time_ns_1_RNIV1DN9_0_21_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire elapsed_time_ns_1_RNI46CN9_0_17_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire bfn_14_13_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire bfn_14_14_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire delay_hc_input_c_g;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire elapsed_time_ns_1_RNIG23T9_0_4_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire elapsed_time_ns_1_RNI13CN9_0_14_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire elapsed_time_ns_1_RNI25DN9_0_24_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire bfn_15_10_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_15_11_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_15_12_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire bfn_15_13_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.N_163_i_g ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire bfn_15_17_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_15_18_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire bfn_15_19_0_;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire bfn_15_20_0_;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_15_21_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire bfn_15_22_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire bfn_15_23_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire bfn_15_24_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_29 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_27 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_31 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire elapsed_time_ns_1_RNI35CN9_0_16_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire bfn_16_13_0_;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire bfn_16_14_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire bfn_16_15_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_4 ;
    wire \current_shift_inst.un38_control_input_0_s1_5 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_0_s1_3 ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_28 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire bfn_17_3_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_17_4_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire bfn_17_5_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_17_6_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_165_i ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_17_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_17_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_17_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_166_i ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_17_11_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_17_12_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_17_13_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_17_14_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire bfn_17_15_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ;
    wire \current_shift_inst.un38_control_input_0_s0_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ;
    wire \current_shift_inst.un38_control_input_0_s0_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire bfn_17_16_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire bfn_17_17_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.N_1619_i ;
    wire \current_shift_inst.control_input_1 ;
    wire bfn_17_19_0_;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_17_20_0_;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_axb_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_axb_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.control_input_cry_13 ;
    wire \current_shift_inst.control_input_axb_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire \current_shift_inst.control_input_cry_14 ;
    wire \current_shift_inst.control_input_cry_15 ;
    wire \current_shift_inst.control_input_axb_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire bfn_17_21_0_;
    wire \current_shift_inst.control_input_axb_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.control_input_cry_16 ;
    wire \current_shift_inst.control_input_axb_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.control_input_cry_17 ;
    wire \current_shift_inst.control_input_axb_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.control_input_cry_18 ;
    wire \current_shift_inst.control_input_axb_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.control_input_cry_19 ;
    wire \current_shift_inst.control_input_axb_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.control_input_cry_20 ;
    wire \current_shift_inst.control_input_axb_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.control_input_cry_21 ;
    wire \current_shift_inst.control_input_axb_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.control_input_cry_22 ;
    wire \current_shift_inst.control_input_cry_23 ;
    wire \current_shift_inst.control_input_axb_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire bfn_17_22_0_;
    wire \current_shift_inst.control_input_axb_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.control_input_cry_24 ;
    wire \current_shift_inst.control_input_axb_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ;
    wire \current_shift_inst.control_input_cry_25 ;
    wire \current_shift_inst.control_input_axb_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ;
    wire \current_shift_inst.control_input_cry_26 ;
    wire \current_shift_inst.control_input_axb_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ;
    wire \current_shift_inst.control_input_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ;
    wire \current_shift_inst.control_input_cry_28 ;
    wire \current_shift_inst.control_input_cry_29 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.control_input_axb_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire bfn_17_23_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire bfn_17_24_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire bfn_17_25_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire bfn_17_26_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_47_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_46_21 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \current_shift_inst.timer_s1.N_164_i ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ;
    wire state_3;
    wire s1_phy_c;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_163_i ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire bfn_18_23_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire bfn_18_24_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire bfn_18_25_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire bfn_18_26_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.N_77_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.N_46_16 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire pwm_duty_input_9;
    wire \current_shift_inst.PI_CTRL.N_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ;
    wire pwm_duty_input_10;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire pwm_duty_input_7;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire pwm_duty_input_6;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire pwm_duty_input_5;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire pwm_duty_input_8;
    wire pwm_duty_input_3;
    wire pwm_duty_input_0;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire pwm_duty_input_1;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.N_97_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire \current_shift_inst.PI_CTRL.N_120 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_98_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__23306),
            .RESETB(N__35876),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42212),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42345),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__40358,N__40283,N__43367,N__40259,N__40481,N__40454,N__43391,N__43346,N__43502,N__40310,N__40337,N__40235,N__43475,N__40160,N__43325,N__43442}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__42347,dangling_wire_45,N__42346}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42704),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42761),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__52734,N__52737,N__52735,N__52738,N__52736,N__52853,N__52970,N__52667,N__53063,N__53009,N__52952,N__52964,N__52913,N__52934,N__52958}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,N__42763,dangling_wire_108,N__42762}),
            .OHOLDTOP(),
            .O({dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_0_14 ,\pwm_generator_inst.O_0_13 ,\pwm_generator_inst.O_0_12 ,\pwm_generator_inst.O_0_11 ,\pwm_generator_inst.O_0_10 ,\pwm_generator_inst.O_0_9 ,\pwm_generator_inst.O_0_8 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_0_6 ,\pwm_generator_inst.O_0_5 ,\pwm_generator_inst.O_0_4 ,\pwm_generator_inst.O_0_3 ,\pwm_generator_inst.O_0_2 ,\pwm_generator_inst.O_0_1 ,\pwm_generator_inst.O_0_0 }));
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42489),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42480),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136}),
            .ADDSUBBOT(),
            .A({dangling_wire_137,N__22769,N__22805,N__22844,N__29846,N__21662,N__21746,N__21701,N__21722,N__21683,N__21788,N__21767,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141}),
            .C({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157}),
            .B({dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,N__42481,N__42488,N__42484,N__42487,N__42482,dangling_wire_164,dangling_wire_165,N__42486,N__42483,N__42485}),
            .OHOLDTOP(),
            .O({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,\pwm_generator_inst.un5_threshold_1_26 ,\pwm_generator_inst.un5_threshold_1_25 ,\pwm_generator_inst.un5_threshold_1_24 ,\pwm_generator_inst.un5_threshold_1_23 ,\pwm_generator_inst.un5_threshold_1_22 ,\pwm_generator_inst.un5_threshold_1_21 ,\pwm_generator_inst.un5_threshold_1_20 ,\pwm_generator_inst.un5_threshold_1_19 ,\pwm_generator_inst.un5_threshold_1_18 ,\pwm_generator_inst.un5_threshold_1_17 ,\pwm_generator_inst.un5_threshold_1_16 ,\pwm_generator_inst.un5_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.O_11 ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42091),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42097),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186}),
            .ADDSUBBOT(),
            .A({N__52796,N__52788,N__52795,N__52787,N__52794,N__52786,N__52793,N__52785,N__52791,N__52783,N__52790,N__52784,N__52792,N__52782,N__52789,N__52781}),
            .C({dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202}),
            .B({dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,N__42099,dangling_wire_216,N__42098}),
            .OHOLDTOP(),
            .O({dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42019),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__41996),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251}),
            .ADDSUBBOT(),
            .A({dangling_wire_252,N__23075,N__22874,N__22889,N__22904,N__22919,N__22934,N__22949,N__22964,N__22979,N__22994,N__22619,N__22634,N__22667,N__22703,N__22733}),
            .C({dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268}),
            .B({dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,N__41997,N__42004,N__42000,N__42003,N__41998,dangling_wire_275,dangling_wire_276,N__42002,N__41999,N__42001}),
            .OHOLDTOP(),
            .O({dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,\pwm_generator_inst.un5_threshold_2_1_16 ,\pwm_generator_inst.un5_threshold_2_1_15 ,\pwm_generator_inst.un5_threshold_2_14 ,\pwm_generator_inst.un5_threshold_2_13 ,\pwm_generator_inst.un5_threshold_2_12 ,\pwm_generator_inst.un5_threshold_2_11 ,\pwm_generator_inst.un5_threshold_2_10 ,\pwm_generator_inst.un5_threshold_2_9 ,\pwm_generator_inst.un5_threshold_2_8 ,\pwm_generator_inst.un5_threshold_2_7 ,\pwm_generator_inst.un5_threshold_2_6 ,\pwm_generator_inst.un5_threshold_2_5 ,\pwm_generator_inst.un5_threshold_2_4 ,\pwm_generator_inst.un5_threshold_2_3 ,\pwm_generator_inst.un5_threshold_2_2 ,\pwm_generator_inst.un5_threshold_2_1 ,\pwm_generator_inst.un5_threshold_2_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__42211),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__42605),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .ADDSUBBOT(),
            .A({dangling_wire_308,N__50375,N__43526,N__50309,N__50258,N__50213,N__50357,N__50282,N__48923,N__48965,N__43421,N__48947,N__50333,N__50237,N__48989,N__53891}),
            .C({dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324}),
            .B({dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,N__42607,dangling_wire_338,N__42606}),
            .OHOLDTOP(),
            .O({dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__54405),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__54407),
            .DIN(N__54406),
            .DOUT(N__54405),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__54407),
            .PADOUT(N__54406),
            .PADIN(N__54405),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__54396),
            .DIN(N__54395),
            .DOUT(N__54394),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__54396),
            .PADOUT(N__54395),
            .PADIN(N__54394),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24023),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__54387),
            .DIN(N__54386),
            .DOUT(N__54385),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__54387),
            .PADOUT(N__54386),
            .PADIN(N__54385),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__54378),
            .DIN(N__54377),
            .DOUT(N__54376),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__54378),
            .PADOUT(N__54377),
            .PADIN(N__54376),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__49097),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__54369),
            .DIN(N__54368),
            .DOUT(N__54367),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__54369),
            .PADOUT(N__54368),
            .PADIN(N__54367),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26609),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__54360),
            .DIN(N__54359),
            .DOUT(N__54358),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__54360),
            .PADOUT(N__54359),
            .PADIN(N__54358),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__54351),
            .DIN(N__54350),
            .DOUT(N__54349),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__54351),
            .PADOUT(N__54350),
            .PADIN(N__54349),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28670),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__54342),
            .DIN(N__54341),
            .DOUT(N__54340),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__54342),
            .PADOUT(N__54341),
            .PADIN(N__54340),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__54333),
            .DIN(N__54332),
            .DOUT(N__54331),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__54333),
            .PADOUT(N__54332),
            .PADIN(N__54331),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__54324),
            .DIN(N__54323),
            .DOUT(N__54322),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__54324),
            .PADOUT(N__54323),
            .PADIN(N__54322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__54315),
            .DIN(N__54314),
            .DOUT(N__54313),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__54315),
            .PADOUT(N__54314),
            .PADIN(N__54313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__30698),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__54306),
            .DIN(N__54305),
            .DOUT(N__54304),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__54306),
            .PADOUT(N__54305),
            .PADIN(N__54304),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__54297),
            .DIN(N__54296),
            .DOUT(N__54295),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__54297),
            .PADOUT(N__54296),
            .PADIN(N__54295),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__12659 (
            .O(N__54278),
            .I(N__54275));
    InMux I__12658 (
            .O(N__54275),
            .I(N__54269));
    InMux I__12657 (
            .O(N__54274),
            .I(N__54269));
    LocalMux I__12656 (
            .O(N__54269),
            .I(N__54266));
    Odrv4 I__12655 (
            .O(N__54266),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__12654 (
            .O(N__54263),
            .I(N__54252));
    InMux I__12653 (
            .O(N__54262),
            .I(N__54252));
    InMux I__12652 (
            .O(N__54261),
            .I(N__54252));
    CascadeMux I__12651 (
            .O(N__54260),
            .I(N__54249));
    InMux I__12650 (
            .O(N__54259),
            .I(N__54243));
    LocalMux I__12649 (
            .O(N__54252),
            .I(N__54240));
    InMux I__12648 (
            .O(N__54249),
            .I(N__54237));
    InMux I__12647 (
            .O(N__54248),
            .I(N__54232));
    InMux I__12646 (
            .O(N__54247),
            .I(N__54232));
    InMux I__12645 (
            .O(N__54246),
            .I(N__54229));
    LocalMux I__12644 (
            .O(N__54243),
            .I(N__54222));
    Span4Mux_v I__12643 (
            .O(N__54240),
            .I(N__54222));
    LocalMux I__12642 (
            .O(N__54237),
            .I(N__54222));
    LocalMux I__12641 (
            .O(N__54232),
            .I(N__54217));
    LocalMux I__12640 (
            .O(N__54229),
            .I(N__54217));
    Span4Mux_h I__12639 (
            .O(N__54222),
            .I(N__54214));
    Span4Mux_s2_h I__12638 (
            .O(N__54217),
            .I(N__54211));
    Span4Mux_v I__12637 (
            .O(N__54214),
            .I(N__54208));
    Span4Mux_v I__12636 (
            .O(N__54211),
            .I(N__54205));
    Span4Mux_v I__12635 (
            .O(N__54208),
            .I(N__54202));
    Span4Mux_v I__12634 (
            .O(N__54205),
            .I(N__54199));
    Odrv4 I__12633 (
            .O(N__54202),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10 ));
    Odrv4 I__12632 (
            .O(N__54199),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10 ));
    CascadeMux I__12631 (
            .O(N__54194),
            .I(\current_shift_inst.PI_CTRL.N_97_cascade_ ));
    InMux I__12630 (
            .O(N__54191),
            .I(N__54187));
    InMux I__12629 (
            .O(N__54190),
            .I(N__54184));
    LocalMux I__12628 (
            .O(N__54187),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    LocalMux I__12627 (
            .O(N__54184),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    InMux I__12626 (
            .O(N__54179),
            .I(N__54170));
    InMux I__12625 (
            .O(N__54178),
            .I(N__54170));
    InMux I__12624 (
            .O(N__54177),
            .I(N__54170));
    LocalMux I__12623 (
            .O(N__54170),
            .I(\current_shift_inst.PI_CTRL.N_120 ));
    InMux I__12622 (
            .O(N__54167),
            .I(N__54161));
    InMux I__12621 (
            .O(N__54166),
            .I(N__54158));
    InMux I__12620 (
            .O(N__54165),
            .I(N__54155));
    InMux I__12619 (
            .O(N__54164),
            .I(N__54152));
    LocalMux I__12618 (
            .O(N__54161),
            .I(N__54147));
    LocalMux I__12617 (
            .O(N__54158),
            .I(N__54147));
    LocalMux I__12616 (
            .O(N__54155),
            .I(N__54144));
    LocalMux I__12615 (
            .O(N__54152),
            .I(N__54141));
    Span4Mux_v I__12614 (
            .O(N__54147),
            .I(N__54138));
    Span4Mux_v I__12613 (
            .O(N__54144),
            .I(N__54133));
    Span4Mux_s2_h I__12612 (
            .O(N__54141),
            .I(N__54133));
    Span4Mux_v I__12611 (
            .O(N__54138),
            .I(N__54130));
    Span4Mux_v I__12610 (
            .O(N__54133),
            .I(N__54127));
    Span4Mux_h I__12609 (
            .O(N__54130),
            .I(N__54124));
    Span4Mux_h I__12608 (
            .O(N__54127),
            .I(N__54121));
    Odrv4 I__12607 (
            .O(N__54124),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__12606 (
            .O(N__54121),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__12605 (
            .O(N__54116),
            .I(N__54111));
    InMux I__12604 (
            .O(N__54115),
            .I(N__54108));
    InMux I__12603 (
            .O(N__54114),
            .I(N__54105));
    LocalMux I__12602 (
            .O(N__54111),
            .I(N__54098));
    LocalMux I__12601 (
            .O(N__54108),
            .I(N__54098));
    LocalMux I__12600 (
            .O(N__54105),
            .I(N__54098));
    Span12Mux_v I__12599 (
            .O(N__54098),
            .I(N__54095));
    Odrv12 I__12598 (
            .O(N__54095),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__12597 (
            .O(N__54092),
            .I(N__54080));
    InMux I__12596 (
            .O(N__54091),
            .I(N__54080));
    InMux I__12595 (
            .O(N__54090),
            .I(N__54073));
    InMux I__12594 (
            .O(N__54089),
            .I(N__54073));
    InMux I__12593 (
            .O(N__54088),
            .I(N__54073));
    InMux I__12592 (
            .O(N__54087),
            .I(N__54068));
    InMux I__12591 (
            .O(N__54086),
            .I(N__54068));
    InMux I__12590 (
            .O(N__54085),
            .I(N__54064));
    LocalMux I__12589 (
            .O(N__54080),
            .I(N__54056));
    LocalMux I__12588 (
            .O(N__54073),
            .I(N__54056));
    LocalMux I__12587 (
            .O(N__54068),
            .I(N__54056));
    InMux I__12586 (
            .O(N__54067),
            .I(N__54053));
    LocalMux I__12585 (
            .O(N__54064),
            .I(N__54050));
    InMux I__12584 (
            .O(N__54063),
            .I(N__54047));
    Span4Mux_v I__12583 (
            .O(N__54056),
            .I(N__54042));
    LocalMux I__12582 (
            .O(N__54053),
            .I(N__54042));
    Span4Mux_v I__12581 (
            .O(N__54050),
            .I(N__54037));
    LocalMux I__12580 (
            .O(N__54047),
            .I(N__54037));
    Span4Mux_h I__12579 (
            .O(N__54042),
            .I(N__54034));
    Span4Mux_v I__12578 (
            .O(N__54037),
            .I(N__54031));
    Span4Mux_v I__12577 (
            .O(N__54034),
            .I(N__54028));
    Span4Mux_v I__12576 (
            .O(N__54031),
            .I(N__54025));
    Span4Mux_v I__12575 (
            .O(N__54028),
            .I(N__54022));
    Span4Mux_h I__12574 (
            .O(N__54025),
            .I(N__54019));
    Odrv4 I__12573 (
            .O(N__54022),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__12572 (
            .O(N__54019),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__12571 (
            .O(N__54014),
            .I(N__54011));
    LocalMux I__12570 (
            .O(N__54011),
            .I(N__54007));
    InMux I__12569 (
            .O(N__54010),
            .I(N__54004));
    Odrv4 I__12568 (
            .O(N__54007),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__12567 (
            .O(N__54004),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__12566 (
            .O(N__53999),
            .I(\current_shift_inst.PI_CTRL.N_98_cascade_ ));
    CascadeMux I__12565 (
            .O(N__53996),
            .I(N__53989));
    CascadeMux I__12564 (
            .O(N__53995),
            .I(N__53986));
    CascadeMux I__12563 (
            .O(N__53994),
            .I(N__53983));
    InMux I__12562 (
            .O(N__53993),
            .I(N__53979));
    InMux I__12561 (
            .O(N__53992),
            .I(N__53976));
    InMux I__12560 (
            .O(N__53989),
            .I(N__53973));
    InMux I__12559 (
            .O(N__53986),
            .I(N__53966));
    InMux I__12558 (
            .O(N__53983),
            .I(N__53966));
    InMux I__12557 (
            .O(N__53982),
            .I(N__53966));
    LocalMux I__12556 (
            .O(N__53979),
            .I(N__53960));
    LocalMux I__12555 (
            .O(N__53976),
            .I(N__53960));
    LocalMux I__12554 (
            .O(N__53973),
            .I(N__53957));
    LocalMux I__12553 (
            .O(N__53966),
            .I(N__53954));
    InMux I__12552 (
            .O(N__53965),
            .I(N__53951));
    Span4Mux_s2_h I__12551 (
            .O(N__53960),
            .I(N__53948));
    Span4Mux_s2_h I__12550 (
            .O(N__53957),
            .I(N__53943));
    Span4Mux_s2_h I__12549 (
            .O(N__53954),
            .I(N__53943));
    LocalMux I__12548 (
            .O(N__53951),
            .I(N__53940));
    Span4Mux_v I__12547 (
            .O(N__53948),
            .I(N__53937));
    Span4Mux_v I__12546 (
            .O(N__53943),
            .I(N__53934));
    Span4Mux_s2_h I__12545 (
            .O(N__53940),
            .I(N__53931));
    Span4Mux_v I__12544 (
            .O(N__53937),
            .I(N__53928));
    Span4Mux_v I__12543 (
            .O(N__53934),
            .I(N__53925));
    Span4Mux_v I__12542 (
            .O(N__53931),
            .I(N__53922));
    Odrv4 I__12541 (
            .O(N__53928),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__12540 (
            .O(N__53925),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__12539 (
            .O(N__53922),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__12538 (
            .O(N__53915),
            .I(N__53912));
    LocalMux I__12537 (
            .O(N__53912),
            .I(N__53908));
    InMux I__12536 (
            .O(N__53911),
            .I(N__53905));
    Odrv4 I__12535 (
            .O(N__53908),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    LocalMux I__12534 (
            .O(N__53905),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__12533 (
            .O(N__53900),
            .I(N__53897));
    LocalMux I__12532 (
            .O(N__53897),
            .I(N__53894));
    Odrv12 I__12531 (
            .O(N__53894),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__12530 (
            .O(N__53891),
            .I(N__53887));
    InMux I__12529 (
            .O(N__53890),
            .I(N__53884));
    LocalMux I__12528 (
            .O(N__53887),
            .I(N__53881));
    LocalMux I__12527 (
            .O(N__53884),
            .I(N__53878));
    Span4Mux_v I__12526 (
            .O(N__53881),
            .I(N__53875));
    Span4Mux_h I__12525 (
            .O(N__53878),
            .I(N__53872));
    Span4Mux_h I__12524 (
            .O(N__53875),
            .I(N__53869));
    Span4Mux_h I__12523 (
            .O(N__53872),
            .I(N__53864));
    Span4Mux_h I__12522 (
            .O(N__53869),
            .I(N__53864));
    Odrv4 I__12521 (
            .O(N__53864),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__12520 (
            .O(N__53861),
            .I(N__53858));
    LocalMux I__12519 (
            .O(N__53858),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    ClkMux I__12518 (
            .O(N__53855),
            .I(N__53468));
    ClkMux I__12517 (
            .O(N__53854),
            .I(N__53468));
    ClkMux I__12516 (
            .O(N__53853),
            .I(N__53468));
    ClkMux I__12515 (
            .O(N__53852),
            .I(N__53468));
    ClkMux I__12514 (
            .O(N__53851),
            .I(N__53468));
    ClkMux I__12513 (
            .O(N__53850),
            .I(N__53468));
    ClkMux I__12512 (
            .O(N__53849),
            .I(N__53468));
    ClkMux I__12511 (
            .O(N__53848),
            .I(N__53468));
    ClkMux I__12510 (
            .O(N__53847),
            .I(N__53468));
    ClkMux I__12509 (
            .O(N__53846),
            .I(N__53468));
    ClkMux I__12508 (
            .O(N__53845),
            .I(N__53468));
    ClkMux I__12507 (
            .O(N__53844),
            .I(N__53468));
    ClkMux I__12506 (
            .O(N__53843),
            .I(N__53468));
    ClkMux I__12505 (
            .O(N__53842),
            .I(N__53468));
    ClkMux I__12504 (
            .O(N__53841),
            .I(N__53468));
    ClkMux I__12503 (
            .O(N__53840),
            .I(N__53468));
    ClkMux I__12502 (
            .O(N__53839),
            .I(N__53468));
    ClkMux I__12501 (
            .O(N__53838),
            .I(N__53468));
    ClkMux I__12500 (
            .O(N__53837),
            .I(N__53468));
    ClkMux I__12499 (
            .O(N__53836),
            .I(N__53468));
    ClkMux I__12498 (
            .O(N__53835),
            .I(N__53468));
    ClkMux I__12497 (
            .O(N__53834),
            .I(N__53468));
    ClkMux I__12496 (
            .O(N__53833),
            .I(N__53468));
    ClkMux I__12495 (
            .O(N__53832),
            .I(N__53468));
    ClkMux I__12494 (
            .O(N__53831),
            .I(N__53468));
    ClkMux I__12493 (
            .O(N__53830),
            .I(N__53468));
    ClkMux I__12492 (
            .O(N__53829),
            .I(N__53468));
    ClkMux I__12491 (
            .O(N__53828),
            .I(N__53468));
    ClkMux I__12490 (
            .O(N__53827),
            .I(N__53468));
    ClkMux I__12489 (
            .O(N__53826),
            .I(N__53468));
    ClkMux I__12488 (
            .O(N__53825),
            .I(N__53468));
    ClkMux I__12487 (
            .O(N__53824),
            .I(N__53468));
    ClkMux I__12486 (
            .O(N__53823),
            .I(N__53468));
    ClkMux I__12485 (
            .O(N__53822),
            .I(N__53468));
    ClkMux I__12484 (
            .O(N__53821),
            .I(N__53468));
    ClkMux I__12483 (
            .O(N__53820),
            .I(N__53468));
    ClkMux I__12482 (
            .O(N__53819),
            .I(N__53468));
    ClkMux I__12481 (
            .O(N__53818),
            .I(N__53468));
    ClkMux I__12480 (
            .O(N__53817),
            .I(N__53468));
    ClkMux I__12479 (
            .O(N__53816),
            .I(N__53468));
    ClkMux I__12478 (
            .O(N__53815),
            .I(N__53468));
    ClkMux I__12477 (
            .O(N__53814),
            .I(N__53468));
    ClkMux I__12476 (
            .O(N__53813),
            .I(N__53468));
    ClkMux I__12475 (
            .O(N__53812),
            .I(N__53468));
    ClkMux I__12474 (
            .O(N__53811),
            .I(N__53468));
    ClkMux I__12473 (
            .O(N__53810),
            .I(N__53468));
    ClkMux I__12472 (
            .O(N__53809),
            .I(N__53468));
    ClkMux I__12471 (
            .O(N__53808),
            .I(N__53468));
    ClkMux I__12470 (
            .O(N__53807),
            .I(N__53468));
    ClkMux I__12469 (
            .O(N__53806),
            .I(N__53468));
    ClkMux I__12468 (
            .O(N__53805),
            .I(N__53468));
    ClkMux I__12467 (
            .O(N__53804),
            .I(N__53468));
    ClkMux I__12466 (
            .O(N__53803),
            .I(N__53468));
    ClkMux I__12465 (
            .O(N__53802),
            .I(N__53468));
    ClkMux I__12464 (
            .O(N__53801),
            .I(N__53468));
    ClkMux I__12463 (
            .O(N__53800),
            .I(N__53468));
    ClkMux I__12462 (
            .O(N__53799),
            .I(N__53468));
    ClkMux I__12461 (
            .O(N__53798),
            .I(N__53468));
    ClkMux I__12460 (
            .O(N__53797),
            .I(N__53468));
    ClkMux I__12459 (
            .O(N__53796),
            .I(N__53468));
    ClkMux I__12458 (
            .O(N__53795),
            .I(N__53468));
    ClkMux I__12457 (
            .O(N__53794),
            .I(N__53468));
    ClkMux I__12456 (
            .O(N__53793),
            .I(N__53468));
    ClkMux I__12455 (
            .O(N__53792),
            .I(N__53468));
    ClkMux I__12454 (
            .O(N__53791),
            .I(N__53468));
    ClkMux I__12453 (
            .O(N__53790),
            .I(N__53468));
    ClkMux I__12452 (
            .O(N__53789),
            .I(N__53468));
    ClkMux I__12451 (
            .O(N__53788),
            .I(N__53468));
    ClkMux I__12450 (
            .O(N__53787),
            .I(N__53468));
    ClkMux I__12449 (
            .O(N__53786),
            .I(N__53468));
    ClkMux I__12448 (
            .O(N__53785),
            .I(N__53468));
    ClkMux I__12447 (
            .O(N__53784),
            .I(N__53468));
    ClkMux I__12446 (
            .O(N__53783),
            .I(N__53468));
    ClkMux I__12445 (
            .O(N__53782),
            .I(N__53468));
    ClkMux I__12444 (
            .O(N__53781),
            .I(N__53468));
    ClkMux I__12443 (
            .O(N__53780),
            .I(N__53468));
    ClkMux I__12442 (
            .O(N__53779),
            .I(N__53468));
    ClkMux I__12441 (
            .O(N__53778),
            .I(N__53468));
    ClkMux I__12440 (
            .O(N__53777),
            .I(N__53468));
    ClkMux I__12439 (
            .O(N__53776),
            .I(N__53468));
    ClkMux I__12438 (
            .O(N__53775),
            .I(N__53468));
    ClkMux I__12437 (
            .O(N__53774),
            .I(N__53468));
    ClkMux I__12436 (
            .O(N__53773),
            .I(N__53468));
    ClkMux I__12435 (
            .O(N__53772),
            .I(N__53468));
    ClkMux I__12434 (
            .O(N__53771),
            .I(N__53468));
    ClkMux I__12433 (
            .O(N__53770),
            .I(N__53468));
    ClkMux I__12432 (
            .O(N__53769),
            .I(N__53468));
    ClkMux I__12431 (
            .O(N__53768),
            .I(N__53468));
    ClkMux I__12430 (
            .O(N__53767),
            .I(N__53468));
    ClkMux I__12429 (
            .O(N__53766),
            .I(N__53468));
    ClkMux I__12428 (
            .O(N__53765),
            .I(N__53468));
    ClkMux I__12427 (
            .O(N__53764),
            .I(N__53468));
    ClkMux I__12426 (
            .O(N__53763),
            .I(N__53468));
    ClkMux I__12425 (
            .O(N__53762),
            .I(N__53468));
    ClkMux I__12424 (
            .O(N__53761),
            .I(N__53468));
    ClkMux I__12423 (
            .O(N__53760),
            .I(N__53468));
    ClkMux I__12422 (
            .O(N__53759),
            .I(N__53468));
    ClkMux I__12421 (
            .O(N__53758),
            .I(N__53468));
    ClkMux I__12420 (
            .O(N__53757),
            .I(N__53468));
    ClkMux I__12419 (
            .O(N__53756),
            .I(N__53468));
    ClkMux I__12418 (
            .O(N__53755),
            .I(N__53468));
    ClkMux I__12417 (
            .O(N__53754),
            .I(N__53468));
    ClkMux I__12416 (
            .O(N__53753),
            .I(N__53468));
    ClkMux I__12415 (
            .O(N__53752),
            .I(N__53468));
    ClkMux I__12414 (
            .O(N__53751),
            .I(N__53468));
    ClkMux I__12413 (
            .O(N__53750),
            .I(N__53468));
    ClkMux I__12412 (
            .O(N__53749),
            .I(N__53468));
    ClkMux I__12411 (
            .O(N__53748),
            .I(N__53468));
    ClkMux I__12410 (
            .O(N__53747),
            .I(N__53468));
    ClkMux I__12409 (
            .O(N__53746),
            .I(N__53468));
    ClkMux I__12408 (
            .O(N__53745),
            .I(N__53468));
    ClkMux I__12407 (
            .O(N__53744),
            .I(N__53468));
    ClkMux I__12406 (
            .O(N__53743),
            .I(N__53468));
    ClkMux I__12405 (
            .O(N__53742),
            .I(N__53468));
    ClkMux I__12404 (
            .O(N__53741),
            .I(N__53468));
    ClkMux I__12403 (
            .O(N__53740),
            .I(N__53468));
    ClkMux I__12402 (
            .O(N__53739),
            .I(N__53468));
    ClkMux I__12401 (
            .O(N__53738),
            .I(N__53468));
    ClkMux I__12400 (
            .O(N__53737),
            .I(N__53468));
    ClkMux I__12399 (
            .O(N__53736),
            .I(N__53468));
    ClkMux I__12398 (
            .O(N__53735),
            .I(N__53468));
    ClkMux I__12397 (
            .O(N__53734),
            .I(N__53468));
    ClkMux I__12396 (
            .O(N__53733),
            .I(N__53468));
    ClkMux I__12395 (
            .O(N__53732),
            .I(N__53468));
    ClkMux I__12394 (
            .O(N__53731),
            .I(N__53468));
    ClkMux I__12393 (
            .O(N__53730),
            .I(N__53468));
    ClkMux I__12392 (
            .O(N__53729),
            .I(N__53468));
    ClkMux I__12391 (
            .O(N__53728),
            .I(N__53468));
    ClkMux I__12390 (
            .O(N__53727),
            .I(N__53468));
    GlobalMux I__12389 (
            .O(N__53468),
            .I(clk_100mhz_0));
    InMux I__12388 (
            .O(N__53465),
            .I(N__53455));
    InMux I__12387 (
            .O(N__53464),
            .I(N__53452));
    InMux I__12386 (
            .O(N__53463),
            .I(N__53449));
    InMux I__12385 (
            .O(N__53462),
            .I(N__53446));
    InMux I__12384 (
            .O(N__53461),
            .I(N__53443));
    InMux I__12383 (
            .O(N__53460),
            .I(N__53440));
    InMux I__12382 (
            .O(N__53459),
            .I(N__53437));
    InMux I__12381 (
            .O(N__53458),
            .I(N__53434));
    LocalMux I__12380 (
            .O(N__53455),
            .I(N__53431));
    LocalMux I__12379 (
            .O(N__53452),
            .I(N__53428));
    LocalMux I__12378 (
            .O(N__53449),
            .I(N__53425));
    LocalMux I__12377 (
            .O(N__53446),
            .I(N__53419));
    LocalMux I__12376 (
            .O(N__53443),
            .I(N__53397));
    LocalMux I__12375 (
            .O(N__53440),
            .I(N__53359));
    LocalMux I__12374 (
            .O(N__53437),
            .I(N__53351));
    LocalMux I__12373 (
            .O(N__53434),
            .I(N__53332));
    Glb2LocalMux I__12372 (
            .O(N__53431),
            .I(N__53099));
    Glb2LocalMux I__12371 (
            .O(N__53428),
            .I(N__53099));
    Glb2LocalMux I__12370 (
            .O(N__53425),
            .I(N__53099));
    SRMux I__12369 (
            .O(N__53424),
            .I(N__53099));
    SRMux I__12368 (
            .O(N__53423),
            .I(N__53099));
    SRMux I__12367 (
            .O(N__53422),
            .I(N__53099));
    Glb2LocalMux I__12366 (
            .O(N__53419),
            .I(N__53099));
    SRMux I__12365 (
            .O(N__53418),
            .I(N__53099));
    SRMux I__12364 (
            .O(N__53417),
            .I(N__53099));
    SRMux I__12363 (
            .O(N__53416),
            .I(N__53099));
    SRMux I__12362 (
            .O(N__53415),
            .I(N__53099));
    SRMux I__12361 (
            .O(N__53414),
            .I(N__53099));
    SRMux I__12360 (
            .O(N__53413),
            .I(N__53099));
    SRMux I__12359 (
            .O(N__53412),
            .I(N__53099));
    SRMux I__12358 (
            .O(N__53411),
            .I(N__53099));
    SRMux I__12357 (
            .O(N__53410),
            .I(N__53099));
    SRMux I__12356 (
            .O(N__53409),
            .I(N__53099));
    SRMux I__12355 (
            .O(N__53408),
            .I(N__53099));
    SRMux I__12354 (
            .O(N__53407),
            .I(N__53099));
    SRMux I__12353 (
            .O(N__53406),
            .I(N__53099));
    SRMux I__12352 (
            .O(N__53405),
            .I(N__53099));
    SRMux I__12351 (
            .O(N__53404),
            .I(N__53099));
    SRMux I__12350 (
            .O(N__53403),
            .I(N__53099));
    SRMux I__12349 (
            .O(N__53402),
            .I(N__53099));
    SRMux I__12348 (
            .O(N__53401),
            .I(N__53099));
    SRMux I__12347 (
            .O(N__53400),
            .I(N__53099));
    Glb2LocalMux I__12346 (
            .O(N__53397),
            .I(N__53099));
    SRMux I__12345 (
            .O(N__53396),
            .I(N__53099));
    SRMux I__12344 (
            .O(N__53395),
            .I(N__53099));
    SRMux I__12343 (
            .O(N__53394),
            .I(N__53099));
    SRMux I__12342 (
            .O(N__53393),
            .I(N__53099));
    SRMux I__12341 (
            .O(N__53392),
            .I(N__53099));
    SRMux I__12340 (
            .O(N__53391),
            .I(N__53099));
    SRMux I__12339 (
            .O(N__53390),
            .I(N__53099));
    SRMux I__12338 (
            .O(N__53389),
            .I(N__53099));
    SRMux I__12337 (
            .O(N__53388),
            .I(N__53099));
    SRMux I__12336 (
            .O(N__53387),
            .I(N__53099));
    SRMux I__12335 (
            .O(N__53386),
            .I(N__53099));
    SRMux I__12334 (
            .O(N__53385),
            .I(N__53099));
    SRMux I__12333 (
            .O(N__53384),
            .I(N__53099));
    SRMux I__12332 (
            .O(N__53383),
            .I(N__53099));
    SRMux I__12331 (
            .O(N__53382),
            .I(N__53099));
    SRMux I__12330 (
            .O(N__53381),
            .I(N__53099));
    SRMux I__12329 (
            .O(N__53380),
            .I(N__53099));
    SRMux I__12328 (
            .O(N__53379),
            .I(N__53099));
    SRMux I__12327 (
            .O(N__53378),
            .I(N__53099));
    SRMux I__12326 (
            .O(N__53377),
            .I(N__53099));
    SRMux I__12325 (
            .O(N__53376),
            .I(N__53099));
    SRMux I__12324 (
            .O(N__53375),
            .I(N__53099));
    SRMux I__12323 (
            .O(N__53374),
            .I(N__53099));
    SRMux I__12322 (
            .O(N__53373),
            .I(N__53099));
    SRMux I__12321 (
            .O(N__53372),
            .I(N__53099));
    SRMux I__12320 (
            .O(N__53371),
            .I(N__53099));
    SRMux I__12319 (
            .O(N__53370),
            .I(N__53099));
    SRMux I__12318 (
            .O(N__53369),
            .I(N__53099));
    SRMux I__12317 (
            .O(N__53368),
            .I(N__53099));
    SRMux I__12316 (
            .O(N__53367),
            .I(N__53099));
    SRMux I__12315 (
            .O(N__53366),
            .I(N__53099));
    SRMux I__12314 (
            .O(N__53365),
            .I(N__53099));
    SRMux I__12313 (
            .O(N__53364),
            .I(N__53099));
    SRMux I__12312 (
            .O(N__53363),
            .I(N__53099));
    SRMux I__12311 (
            .O(N__53362),
            .I(N__53099));
    Glb2LocalMux I__12310 (
            .O(N__53359),
            .I(N__53099));
    SRMux I__12309 (
            .O(N__53358),
            .I(N__53099));
    SRMux I__12308 (
            .O(N__53357),
            .I(N__53099));
    SRMux I__12307 (
            .O(N__53356),
            .I(N__53099));
    SRMux I__12306 (
            .O(N__53355),
            .I(N__53099));
    SRMux I__12305 (
            .O(N__53354),
            .I(N__53099));
    Glb2LocalMux I__12304 (
            .O(N__53351),
            .I(N__53099));
    SRMux I__12303 (
            .O(N__53350),
            .I(N__53099));
    SRMux I__12302 (
            .O(N__53349),
            .I(N__53099));
    SRMux I__12301 (
            .O(N__53348),
            .I(N__53099));
    SRMux I__12300 (
            .O(N__53347),
            .I(N__53099));
    SRMux I__12299 (
            .O(N__53346),
            .I(N__53099));
    SRMux I__12298 (
            .O(N__53345),
            .I(N__53099));
    SRMux I__12297 (
            .O(N__53344),
            .I(N__53099));
    SRMux I__12296 (
            .O(N__53343),
            .I(N__53099));
    SRMux I__12295 (
            .O(N__53342),
            .I(N__53099));
    SRMux I__12294 (
            .O(N__53341),
            .I(N__53099));
    SRMux I__12293 (
            .O(N__53340),
            .I(N__53099));
    SRMux I__12292 (
            .O(N__53339),
            .I(N__53099));
    SRMux I__12291 (
            .O(N__53338),
            .I(N__53099));
    SRMux I__12290 (
            .O(N__53337),
            .I(N__53099));
    SRMux I__12289 (
            .O(N__53336),
            .I(N__53099));
    SRMux I__12288 (
            .O(N__53335),
            .I(N__53099));
    Glb2LocalMux I__12287 (
            .O(N__53332),
            .I(N__53099));
    SRMux I__12286 (
            .O(N__53331),
            .I(N__53099));
    SRMux I__12285 (
            .O(N__53330),
            .I(N__53099));
    SRMux I__12284 (
            .O(N__53329),
            .I(N__53099));
    SRMux I__12283 (
            .O(N__53328),
            .I(N__53099));
    SRMux I__12282 (
            .O(N__53327),
            .I(N__53099));
    SRMux I__12281 (
            .O(N__53326),
            .I(N__53099));
    SRMux I__12280 (
            .O(N__53325),
            .I(N__53099));
    SRMux I__12279 (
            .O(N__53324),
            .I(N__53099));
    SRMux I__12278 (
            .O(N__53323),
            .I(N__53099));
    SRMux I__12277 (
            .O(N__53322),
            .I(N__53099));
    SRMux I__12276 (
            .O(N__53321),
            .I(N__53099));
    SRMux I__12275 (
            .O(N__53320),
            .I(N__53099));
    SRMux I__12274 (
            .O(N__53319),
            .I(N__53099));
    SRMux I__12273 (
            .O(N__53318),
            .I(N__53099));
    SRMux I__12272 (
            .O(N__53317),
            .I(N__53099));
    SRMux I__12271 (
            .O(N__53316),
            .I(N__53099));
    SRMux I__12270 (
            .O(N__53315),
            .I(N__53099));
    SRMux I__12269 (
            .O(N__53314),
            .I(N__53099));
    SRMux I__12268 (
            .O(N__53313),
            .I(N__53099));
    SRMux I__12267 (
            .O(N__53312),
            .I(N__53099));
    GlobalMux I__12266 (
            .O(N__53099),
            .I(N__53096));
    gio2CtrlBuf I__12265 (
            .O(N__53096),
            .I(red_c_g));
    InMux I__12264 (
            .O(N__53093),
            .I(N__53086));
    InMux I__12263 (
            .O(N__53092),
            .I(N__53086));
    InMux I__12262 (
            .O(N__53091),
            .I(N__53083));
    LocalMux I__12261 (
            .O(N__53086),
            .I(N__53080));
    LocalMux I__12260 (
            .O(N__53083),
            .I(N__53077));
    Span4Mux_v I__12259 (
            .O(N__53080),
            .I(N__53074));
    Span12Mux_s7_h I__12258 (
            .O(N__53077),
            .I(N__53071));
    Span4Mux_h I__12257 (
            .O(N__53074),
            .I(N__53068));
    Odrv12 I__12256 (
            .O(N__53071),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__12255 (
            .O(N__53068),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__12254 (
            .O(N__53063),
            .I(N__53060));
    LocalMux I__12253 (
            .O(N__53060),
            .I(pwm_duty_input_6));
    CascadeMux I__12252 (
            .O(N__53057),
            .I(N__53053));
    CascadeMux I__12251 (
            .O(N__53056),
            .I(N__53050));
    InMux I__12250 (
            .O(N__53053),
            .I(N__53047));
    InMux I__12249 (
            .O(N__53050),
            .I(N__53044));
    LocalMux I__12248 (
            .O(N__53047),
            .I(N__53040));
    LocalMux I__12247 (
            .O(N__53044),
            .I(N__53037));
    InMux I__12246 (
            .O(N__53043),
            .I(N__53034));
    Span4Mux_v I__12245 (
            .O(N__53040),
            .I(N__53031));
    Span4Mux_s2_h I__12244 (
            .O(N__53037),
            .I(N__53026));
    LocalMux I__12243 (
            .O(N__53034),
            .I(N__53026));
    Span4Mux_v I__12242 (
            .O(N__53031),
            .I(N__53023));
    Span4Mux_v I__12241 (
            .O(N__53026),
            .I(N__53020));
    Span4Mux_h I__12240 (
            .O(N__53023),
            .I(N__53017));
    Span4Mux_h I__12239 (
            .O(N__53020),
            .I(N__53014));
    Odrv4 I__12238 (
            .O(N__53017),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__12237 (
            .O(N__53014),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__12236 (
            .O(N__53009),
            .I(N__53006));
    LocalMux I__12235 (
            .O(N__53006),
            .I(pwm_duty_input_5));
    InMux I__12234 (
            .O(N__53003),
            .I(N__52999));
    InMux I__12233 (
            .O(N__53002),
            .I(N__52996));
    LocalMux I__12232 (
            .O(N__52999),
            .I(N__52993));
    LocalMux I__12231 (
            .O(N__52996),
            .I(N__52990));
    Span4Mux_v I__12230 (
            .O(N__52993),
            .I(N__52984));
    Span4Mux_v I__12229 (
            .O(N__52990),
            .I(N__52984));
    InMux I__12228 (
            .O(N__52989),
            .I(N__52981));
    Sp12to4 I__12227 (
            .O(N__52984),
            .I(N__52976));
    LocalMux I__12226 (
            .O(N__52981),
            .I(N__52976));
    Span12Mux_s7_h I__12225 (
            .O(N__52976),
            .I(N__52973));
    Odrv12 I__12224 (
            .O(N__52973),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__12223 (
            .O(N__52970),
            .I(N__52967));
    LocalMux I__12222 (
            .O(N__52967),
            .I(pwm_duty_input_8));
    InMux I__12221 (
            .O(N__52964),
            .I(N__52961));
    LocalMux I__12220 (
            .O(N__52961),
            .I(pwm_duty_input_3));
    InMux I__12219 (
            .O(N__52958),
            .I(N__52955));
    LocalMux I__12218 (
            .O(N__52955),
            .I(pwm_duty_input_0));
    InMux I__12217 (
            .O(N__52952),
            .I(N__52949));
    LocalMux I__12216 (
            .O(N__52949),
            .I(pwm_duty_input_4));
    InMux I__12215 (
            .O(N__52946),
            .I(N__52943));
    LocalMux I__12214 (
            .O(N__52943),
            .I(N__52940));
    Span12Mux_s7_h I__12213 (
            .O(N__52940),
            .I(N__52937));
    Odrv12 I__12212 (
            .O(N__52937),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__12211 (
            .O(N__52934),
            .I(N__52931));
    LocalMux I__12210 (
            .O(N__52931),
            .I(pwm_duty_input_1));
    InMux I__12209 (
            .O(N__52928),
            .I(N__52925));
    LocalMux I__12208 (
            .O(N__52925),
            .I(N__52922));
    Sp12to4 I__12207 (
            .O(N__52922),
            .I(N__52919));
    Span12Mux_v I__12206 (
            .O(N__52919),
            .I(N__52916));
    Odrv12 I__12205 (
            .O(N__52916),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__12204 (
            .O(N__52913),
            .I(N__52910));
    LocalMux I__12203 (
            .O(N__52910),
            .I(pwm_duty_input_2));
    InMux I__12202 (
            .O(N__52907),
            .I(N__52904));
    LocalMux I__12201 (
            .O(N__52904),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    InMux I__12200 (
            .O(N__52901),
            .I(N__52898));
    LocalMux I__12199 (
            .O(N__52898),
            .I(N__52895));
    Span4Mux_h I__12198 (
            .O(N__52895),
            .I(N__52892));
    Odrv4 I__12197 (
            .O(N__52892),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__12196 (
            .O(N__52889),
            .I(N__52886));
    LocalMux I__12195 (
            .O(N__52886),
            .I(N__52883));
    Odrv4 I__12194 (
            .O(N__52883),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    CascadeMux I__12193 (
            .O(N__52880),
            .I(N__52877));
    InMux I__12192 (
            .O(N__52877),
            .I(N__52874));
    LocalMux I__12191 (
            .O(N__52874),
            .I(N__52871));
    Span4Mux_v I__12190 (
            .O(N__52871),
            .I(N__52868));
    Odrv4 I__12189 (
            .O(N__52868),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__12188 (
            .O(N__52865),
            .I(N__52862));
    LocalMux I__12187 (
            .O(N__52862),
            .I(N__52859));
    Span4Mux_h I__12186 (
            .O(N__52859),
            .I(N__52856));
    Odrv4 I__12185 (
            .O(N__52856),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__12184 (
            .O(N__52853),
            .I(N__52850));
    LocalMux I__12183 (
            .O(N__52850),
            .I(N__52847));
    Span4Mux_s1_h I__12182 (
            .O(N__52847),
            .I(N__52844));
    Odrv4 I__12181 (
            .O(N__52844),
            .I(pwm_duty_input_9));
    CascadeMux I__12180 (
            .O(N__52841),
            .I(\current_shift_inst.PI_CTRL.N_31_cascade_ ));
    CascadeMux I__12179 (
            .O(N__52838),
            .I(N__52835));
    InMux I__12178 (
            .O(N__52835),
            .I(N__52832));
    LocalMux I__12177 (
            .O(N__52832),
            .I(N__52827));
    InMux I__12176 (
            .O(N__52831),
            .I(N__52824));
    InMux I__12175 (
            .O(N__52830),
            .I(N__52821));
    Span4Mux_v I__12174 (
            .O(N__52827),
            .I(N__52814));
    LocalMux I__12173 (
            .O(N__52824),
            .I(N__52814));
    LocalMux I__12172 (
            .O(N__52821),
            .I(N__52814));
    Span4Mux_v I__12171 (
            .O(N__52814),
            .I(N__52811));
    Span4Mux_h I__12170 (
            .O(N__52811),
            .I(N__52808));
    Odrv4 I__12169 (
            .O(N__52808),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    CascadeMux I__12168 (
            .O(N__52805),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    InMux I__12167 (
            .O(N__52802),
            .I(N__52799));
    LocalMux I__12166 (
            .O(N__52799),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ));
    InMux I__12165 (
            .O(N__52796),
            .I(N__52764));
    InMux I__12164 (
            .O(N__52795),
            .I(N__52764));
    InMux I__12163 (
            .O(N__52794),
            .I(N__52764));
    InMux I__12162 (
            .O(N__52793),
            .I(N__52764));
    InMux I__12161 (
            .O(N__52792),
            .I(N__52764));
    InMux I__12160 (
            .O(N__52791),
            .I(N__52764));
    InMux I__12159 (
            .O(N__52790),
            .I(N__52764));
    InMux I__12158 (
            .O(N__52789),
            .I(N__52764));
    InMux I__12157 (
            .O(N__52788),
            .I(N__52747));
    InMux I__12156 (
            .O(N__52787),
            .I(N__52747));
    InMux I__12155 (
            .O(N__52786),
            .I(N__52747));
    InMux I__12154 (
            .O(N__52785),
            .I(N__52747));
    InMux I__12153 (
            .O(N__52784),
            .I(N__52747));
    InMux I__12152 (
            .O(N__52783),
            .I(N__52747));
    InMux I__12151 (
            .O(N__52782),
            .I(N__52747));
    InMux I__12150 (
            .O(N__52781),
            .I(N__52747));
    LocalMux I__12149 (
            .O(N__52764),
            .I(N__52742));
    LocalMux I__12148 (
            .O(N__52747),
            .I(N__52742));
    Span4Mux_v I__12147 (
            .O(N__52742),
            .I(N__52739));
    Sp12to4 I__12146 (
            .O(N__52739),
            .I(N__52731));
    InMux I__12145 (
            .O(N__52738),
            .I(N__52726));
    InMux I__12144 (
            .O(N__52737),
            .I(N__52726));
    InMux I__12143 (
            .O(N__52736),
            .I(N__52719));
    InMux I__12142 (
            .O(N__52735),
            .I(N__52719));
    InMux I__12141 (
            .O(N__52734),
            .I(N__52719));
    Span12Mux_s8_h I__12140 (
            .O(N__52731),
            .I(N__52716));
    LocalMux I__12139 (
            .O(N__52726),
            .I(N__52711));
    LocalMux I__12138 (
            .O(N__52719),
            .I(N__52711));
    Span12Mux_h I__12137 (
            .O(N__52716),
            .I(N__52708));
    Odrv4 I__12136 (
            .O(N__52711),
            .I(pwm_duty_input_10));
    Odrv12 I__12135 (
            .O(N__52708),
            .I(pwm_duty_input_10));
    InMux I__12134 (
            .O(N__52703),
            .I(N__52700));
    LocalMux I__12133 (
            .O(N__52700),
            .I(N__52695));
    InMux I__12132 (
            .O(N__52699),
            .I(N__52690));
    InMux I__12131 (
            .O(N__52698),
            .I(N__52690));
    Span4Mux_h I__12130 (
            .O(N__52695),
            .I(N__52687));
    LocalMux I__12129 (
            .O(N__52690),
            .I(N__52684));
    Span4Mux_v I__12128 (
            .O(N__52687),
            .I(N__52681));
    Span4Mux_v I__12127 (
            .O(N__52684),
            .I(N__52678));
    Span4Mux_v I__12126 (
            .O(N__52681),
            .I(N__52675));
    Span4Mux_h I__12125 (
            .O(N__52678),
            .I(N__52672));
    Odrv4 I__12124 (
            .O(N__52675),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__12123 (
            .O(N__52672),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__12122 (
            .O(N__52667),
            .I(N__52664));
    LocalMux I__12121 (
            .O(N__52664),
            .I(N__52661));
    Odrv4 I__12120 (
            .O(N__52661),
            .I(pwm_duty_input_7));
    InMux I__12119 (
            .O(N__52658),
            .I(N__52655));
    LocalMux I__12118 (
            .O(N__52655),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    CascadeMux I__12117 (
            .O(N__52652),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    InMux I__12116 (
            .O(N__52649),
            .I(N__52643));
    InMux I__12115 (
            .O(N__52648),
            .I(N__52643));
    LocalMux I__12114 (
            .O(N__52643),
            .I(N__52640));
    Odrv4 I__12113 (
            .O(N__52640),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__12112 (
            .O(N__52637),
            .I(N__52634));
    LocalMux I__12111 (
            .O(N__52634),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__12110 (
            .O(N__52631),
            .I(N__52628));
    LocalMux I__12109 (
            .O(N__52628),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__12108 (
            .O(N__52625),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ));
    InMux I__12107 (
            .O(N__52622),
            .I(N__52618));
    InMux I__12106 (
            .O(N__52621),
            .I(N__52615));
    LocalMux I__12105 (
            .O(N__52618),
            .I(N__52612));
    LocalMux I__12104 (
            .O(N__52615),
            .I(N__52609));
    Span4Mux_h I__12103 (
            .O(N__52612),
            .I(N__52606));
    Odrv4 I__12102 (
            .O(N__52609),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    Odrv4 I__12101 (
            .O(N__52606),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__12100 (
            .O(N__52601),
            .I(N__52597));
    InMux I__12099 (
            .O(N__52600),
            .I(N__52594));
    LocalMux I__12098 (
            .O(N__52597),
            .I(N__52591));
    LocalMux I__12097 (
            .O(N__52594),
            .I(N__52588));
    Span4Mux_h I__12096 (
            .O(N__52591),
            .I(N__52585));
    Odrv4 I__12095 (
            .O(N__52588),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    Odrv4 I__12094 (
            .O(N__52585),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__12093 (
            .O(N__52580),
            .I(N__52576));
    InMux I__12092 (
            .O(N__52579),
            .I(N__52573));
    LocalMux I__12091 (
            .O(N__52576),
            .I(N__52570));
    LocalMux I__12090 (
            .O(N__52573),
            .I(N__52567));
    Span4Mux_h I__12089 (
            .O(N__52570),
            .I(N__52564));
    Odrv4 I__12088 (
            .O(N__52567),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    Odrv4 I__12087 (
            .O(N__52564),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    CascadeMux I__12086 (
            .O(N__52559),
            .I(N__52555));
    InMux I__12085 (
            .O(N__52558),
            .I(N__52550));
    InMux I__12084 (
            .O(N__52555),
            .I(N__52550));
    LocalMux I__12083 (
            .O(N__52550),
            .I(N__52547));
    Odrv4 I__12082 (
            .O(N__52547),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__12081 (
            .O(N__52544),
            .I(N__52538));
    InMux I__12080 (
            .O(N__52543),
            .I(N__52538));
    LocalMux I__12079 (
            .O(N__52538),
            .I(N__52535));
    Odrv4 I__12078 (
            .O(N__52535),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__12077 (
            .O(N__52532),
            .I(N__52526));
    InMux I__12076 (
            .O(N__52531),
            .I(N__52526));
    LocalMux I__12075 (
            .O(N__52526),
            .I(N__52523));
    Odrv4 I__12074 (
            .O(N__52523),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__12073 (
            .O(N__52520),
            .I(N__52514));
    InMux I__12072 (
            .O(N__52519),
            .I(N__52514));
    LocalMux I__12071 (
            .O(N__52514),
            .I(N__52511));
    Odrv4 I__12070 (
            .O(N__52511),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    CascadeMux I__12069 (
            .O(N__52508),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    CascadeMux I__12068 (
            .O(N__52505),
            .I(N__52501));
    InMux I__12067 (
            .O(N__52504),
            .I(N__52498));
    InMux I__12066 (
            .O(N__52501),
            .I(N__52495));
    LocalMux I__12065 (
            .O(N__52498),
            .I(N__52490));
    LocalMux I__12064 (
            .O(N__52495),
            .I(N__52490));
    Span4Mux_h I__12063 (
            .O(N__52490),
            .I(N__52487));
    Odrv4 I__12062 (
            .O(N__52487),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__12061 (
            .O(N__52484),
            .I(N__52481));
    LocalMux I__12060 (
            .O(N__52481),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__12059 (
            .O(N__52478),
            .I(N__52475));
    LocalMux I__12058 (
            .O(N__52475),
            .I(N__52472));
    Span4Mux_h I__12057 (
            .O(N__52472),
            .I(N__52469));
    Odrv4 I__12056 (
            .O(N__52469),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    CascadeMux I__12055 (
            .O(N__52466),
            .I(N__52463));
    InMux I__12054 (
            .O(N__52463),
            .I(N__52459));
    InMux I__12053 (
            .O(N__52462),
            .I(N__52456));
    LocalMux I__12052 (
            .O(N__52459),
            .I(N__52451));
    LocalMux I__12051 (
            .O(N__52456),
            .I(N__52448));
    InMux I__12050 (
            .O(N__52455),
            .I(N__52445));
    InMux I__12049 (
            .O(N__52454),
            .I(N__52442));
    Span4Mux_v I__12048 (
            .O(N__52451),
            .I(N__52439));
    Span4Mux_v I__12047 (
            .O(N__52448),
            .I(N__52432));
    LocalMux I__12046 (
            .O(N__52445),
            .I(N__52432));
    LocalMux I__12045 (
            .O(N__52442),
            .I(N__52432));
    Odrv4 I__12044 (
            .O(N__52439),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__12043 (
            .O(N__52432),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__12042 (
            .O(N__52427),
            .I(N__52413));
    InMux I__12041 (
            .O(N__52426),
            .I(N__52408));
    InMux I__12040 (
            .O(N__52425),
            .I(N__52408));
    InMux I__12039 (
            .O(N__52424),
            .I(N__52405));
    InMux I__12038 (
            .O(N__52423),
            .I(N__52402));
    InMux I__12037 (
            .O(N__52422),
            .I(N__52397));
    InMux I__12036 (
            .O(N__52421),
            .I(N__52394));
    InMux I__12035 (
            .O(N__52420),
            .I(N__52389));
    InMux I__12034 (
            .O(N__52419),
            .I(N__52389));
    CascadeMux I__12033 (
            .O(N__52418),
            .I(N__52384));
    InMux I__12032 (
            .O(N__52417),
            .I(N__52379));
    InMux I__12031 (
            .O(N__52416),
            .I(N__52379));
    LocalMux I__12030 (
            .O(N__52413),
            .I(N__52376));
    LocalMux I__12029 (
            .O(N__52408),
            .I(N__52358));
    LocalMux I__12028 (
            .O(N__52405),
            .I(N__52355));
    LocalMux I__12027 (
            .O(N__52402),
            .I(N__52352));
    InMux I__12026 (
            .O(N__52401),
            .I(N__52347));
    InMux I__12025 (
            .O(N__52400),
            .I(N__52347));
    LocalMux I__12024 (
            .O(N__52397),
            .I(N__52344));
    LocalMux I__12023 (
            .O(N__52394),
            .I(N__52339));
    LocalMux I__12022 (
            .O(N__52389),
            .I(N__52339));
    InMux I__12021 (
            .O(N__52388),
            .I(N__52332));
    InMux I__12020 (
            .O(N__52387),
            .I(N__52332));
    InMux I__12019 (
            .O(N__52384),
            .I(N__52332));
    LocalMux I__12018 (
            .O(N__52379),
            .I(N__52329));
    Span4Mux_v I__12017 (
            .O(N__52376),
            .I(N__52326));
    InMux I__12016 (
            .O(N__52375),
            .I(N__52323));
    InMux I__12015 (
            .O(N__52374),
            .I(N__52320));
    InMux I__12014 (
            .O(N__52373),
            .I(N__52307));
    InMux I__12013 (
            .O(N__52372),
            .I(N__52307));
    InMux I__12012 (
            .O(N__52371),
            .I(N__52307));
    InMux I__12011 (
            .O(N__52370),
            .I(N__52307));
    InMux I__12010 (
            .O(N__52369),
            .I(N__52307));
    InMux I__12009 (
            .O(N__52368),
            .I(N__52307));
    InMux I__12008 (
            .O(N__52367),
            .I(N__52304));
    InMux I__12007 (
            .O(N__52366),
            .I(N__52291));
    InMux I__12006 (
            .O(N__52365),
            .I(N__52291));
    InMux I__12005 (
            .O(N__52364),
            .I(N__52291));
    InMux I__12004 (
            .O(N__52363),
            .I(N__52291));
    InMux I__12003 (
            .O(N__52362),
            .I(N__52291));
    InMux I__12002 (
            .O(N__52361),
            .I(N__52291));
    Span4Mux_h I__12001 (
            .O(N__52358),
            .I(N__52284));
    Span4Mux_h I__12000 (
            .O(N__52355),
            .I(N__52284));
    Span4Mux_h I__11999 (
            .O(N__52352),
            .I(N__52284));
    LocalMux I__11998 (
            .O(N__52347),
            .I(N__52275));
    Span4Mux_h I__11997 (
            .O(N__52344),
            .I(N__52275));
    Span4Mux_v I__11996 (
            .O(N__52339),
            .I(N__52275));
    LocalMux I__11995 (
            .O(N__52332),
            .I(N__52275));
    Span4Mux_h I__11994 (
            .O(N__52329),
            .I(N__52268));
    Span4Mux_h I__11993 (
            .O(N__52326),
            .I(N__52268));
    LocalMux I__11992 (
            .O(N__52323),
            .I(N__52268));
    LocalMux I__11991 (
            .O(N__52320),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__11990 (
            .O(N__52307),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__11989 (
            .O(N__52304),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__11988 (
            .O(N__52291),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__11987 (
            .O(N__52284),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__11986 (
            .O(N__52275),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__11985 (
            .O(N__52268),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__11984 (
            .O(N__52253),
            .I(N__52250));
    LocalMux I__11983 (
            .O(N__52250),
            .I(N__52247));
    Span4Mux_h I__11982 (
            .O(N__52247),
            .I(N__52244));
    Odrv4 I__11981 (
            .O(N__52244),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__11980 (
            .O(N__52241),
            .I(N__52230));
    InMux I__11979 (
            .O(N__52240),
            .I(N__52227));
    InMux I__11978 (
            .O(N__52239),
            .I(N__52224));
    InMux I__11977 (
            .O(N__52238),
            .I(N__52216));
    InMux I__11976 (
            .O(N__52237),
            .I(N__52216));
    InMux I__11975 (
            .O(N__52236),
            .I(N__52201));
    InMux I__11974 (
            .O(N__52235),
            .I(N__52198));
    InMux I__11973 (
            .O(N__52234),
            .I(N__52191));
    InMux I__11972 (
            .O(N__52233),
            .I(N__52191));
    LocalMux I__11971 (
            .O(N__52230),
            .I(N__52184));
    LocalMux I__11970 (
            .O(N__52227),
            .I(N__52181));
    LocalMux I__11969 (
            .O(N__52224),
            .I(N__52178));
    InMux I__11968 (
            .O(N__52223),
            .I(N__52173));
    InMux I__11967 (
            .O(N__52222),
            .I(N__52173));
    CEMux I__11966 (
            .O(N__52221),
            .I(N__52170));
    LocalMux I__11965 (
            .O(N__52216),
            .I(N__52167));
    InMux I__11964 (
            .O(N__52215),
            .I(N__52154));
    InMux I__11963 (
            .O(N__52214),
            .I(N__52154));
    InMux I__11962 (
            .O(N__52213),
            .I(N__52154));
    InMux I__11961 (
            .O(N__52212),
            .I(N__52154));
    InMux I__11960 (
            .O(N__52211),
            .I(N__52154));
    InMux I__11959 (
            .O(N__52210),
            .I(N__52154));
    InMux I__11958 (
            .O(N__52209),
            .I(N__52141));
    InMux I__11957 (
            .O(N__52208),
            .I(N__52141));
    InMux I__11956 (
            .O(N__52207),
            .I(N__52141));
    InMux I__11955 (
            .O(N__52206),
            .I(N__52141));
    InMux I__11954 (
            .O(N__52205),
            .I(N__52141));
    InMux I__11953 (
            .O(N__52204),
            .I(N__52141));
    LocalMux I__11952 (
            .O(N__52201),
            .I(N__52136));
    LocalMux I__11951 (
            .O(N__52198),
            .I(N__52136));
    InMux I__11950 (
            .O(N__52197),
            .I(N__52131));
    InMux I__11949 (
            .O(N__52196),
            .I(N__52131));
    LocalMux I__11948 (
            .O(N__52191),
            .I(N__52128));
    InMux I__11947 (
            .O(N__52190),
            .I(N__52125));
    InMux I__11946 (
            .O(N__52189),
            .I(N__52122));
    InMux I__11945 (
            .O(N__52188),
            .I(N__52117));
    InMux I__11944 (
            .O(N__52187),
            .I(N__52117));
    Span4Mux_h I__11943 (
            .O(N__52184),
            .I(N__52112));
    Span4Mux_h I__11942 (
            .O(N__52181),
            .I(N__52112));
    Span4Mux_v I__11941 (
            .O(N__52178),
            .I(N__52109));
    LocalMux I__11940 (
            .O(N__52173),
            .I(N__52106));
    LocalMux I__11939 (
            .O(N__52170),
            .I(N__52095));
    Span4Mux_v I__11938 (
            .O(N__52167),
            .I(N__52095));
    LocalMux I__11937 (
            .O(N__52154),
            .I(N__52095));
    LocalMux I__11936 (
            .O(N__52141),
            .I(N__52095));
    Span4Mux_v I__11935 (
            .O(N__52136),
            .I(N__52095));
    LocalMux I__11934 (
            .O(N__52131),
            .I(N__52090));
    Span12Mux_v I__11933 (
            .O(N__52128),
            .I(N__52090));
    LocalMux I__11932 (
            .O(N__52125),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__11931 (
            .O(N__52122),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__11930 (
            .O(N__52117),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__11929 (
            .O(N__52112),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__11928 (
            .O(N__52109),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv12 I__11927 (
            .O(N__52106),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__11926 (
            .O(N__52095),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv12 I__11925 (
            .O(N__52090),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    CascadeMux I__11924 (
            .O(N__52073),
            .I(N__52069));
    CascadeMux I__11923 (
            .O(N__52072),
            .I(N__52065));
    InMux I__11922 (
            .O(N__52069),
            .I(N__52062));
    InMux I__11921 (
            .O(N__52068),
            .I(N__52059));
    InMux I__11920 (
            .O(N__52065),
            .I(N__52055));
    LocalMux I__11919 (
            .O(N__52062),
            .I(N__52050));
    LocalMux I__11918 (
            .O(N__52059),
            .I(N__52050));
    InMux I__11917 (
            .O(N__52058),
            .I(N__52047));
    LocalMux I__11916 (
            .O(N__52055),
            .I(N__52044));
    Span4Mux_v I__11915 (
            .O(N__52050),
            .I(N__52039));
    LocalMux I__11914 (
            .O(N__52047),
            .I(N__52039));
    Span4Mux_v I__11913 (
            .O(N__52044),
            .I(N__52036));
    Span4Mux_s3_v I__11912 (
            .O(N__52039),
            .I(N__52033));
    Span4Mux_h I__11911 (
            .O(N__52036),
            .I(N__52030));
    Span4Mux_h I__11910 (
            .O(N__52033),
            .I(N__52027));
    Odrv4 I__11909 (
            .O(N__52030),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__11908 (
            .O(N__52027),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__11907 (
            .O(N__52022),
            .I(N__52016));
    InMux I__11906 (
            .O(N__52021),
            .I(N__52016));
    LocalMux I__11905 (
            .O(N__52016),
            .I(N__52013));
    Odrv4 I__11904 (
            .O(N__52013),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    CascadeMux I__11903 (
            .O(N__52010),
            .I(N__52006));
    InMux I__11902 (
            .O(N__52009),
            .I(N__52003));
    InMux I__11901 (
            .O(N__52006),
            .I(N__52000));
    LocalMux I__11900 (
            .O(N__52003),
            .I(N__51995));
    LocalMux I__11899 (
            .O(N__52000),
            .I(N__51995));
    Span4Mux_h I__11898 (
            .O(N__51995),
            .I(N__51992));
    Odrv4 I__11897 (
            .O(N__51992),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    CascadeMux I__11896 (
            .O(N__51989),
            .I(N__51986));
    InMux I__11895 (
            .O(N__51986),
            .I(N__51980));
    InMux I__11894 (
            .O(N__51985),
            .I(N__51980));
    LocalMux I__11893 (
            .O(N__51980),
            .I(N__51977));
    Odrv12 I__11892 (
            .O(N__51977),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__11891 (
            .O(N__51974),
            .I(N__51968));
    InMux I__11890 (
            .O(N__51973),
            .I(N__51968));
    LocalMux I__11889 (
            .O(N__51968),
            .I(N__51965));
    Odrv4 I__11888 (
            .O(N__51965),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    CascadeMux I__11887 (
            .O(N__51962),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ));
    InMux I__11886 (
            .O(N__51959),
            .I(N__51956));
    LocalMux I__11885 (
            .O(N__51956),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    InMux I__11884 (
            .O(N__51953),
            .I(N__51950));
    LocalMux I__11883 (
            .O(N__51950),
            .I(N__51946));
    InMux I__11882 (
            .O(N__51949),
            .I(N__51943));
    Span4Mux_v I__11881 (
            .O(N__51946),
            .I(N__51938));
    LocalMux I__11880 (
            .O(N__51943),
            .I(N__51938));
    Odrv4 I__11879 (
            .O(N__51938),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    CascadeMux I__11878 (
            .O(N__51935),
            .I(N__51932));
    InMux I__11877 (
            .O(N__51932),
            .I(N__51929));
    LocalMux I__11876 (
            .O(N__51929),
            .I(N__51925));
    InMux I__11875 (
            .O(N__51928),
            .I(N__51922));
    Span4Mux_h I__11874 (
            .O(N__51925),
            .I(N__51919));
    LocalMux I__11873 (
            .O(N__51922),
            .I(N__51916));
    Odrv4 I__11872 (
            .O(N__51919),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    Odrv4 I__11871 (
            .O(N__51916),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    CascadeMux I__11870 (
            .O(N__51911),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    InMux I__11869 (
            .O(N__51908),
            .I(N__51902));
    InMux I__11868 (
            .O(N__51907),
            .I(N__51902));
    LocalMux I__11867 (
            .O(N__51902),
            .I(N__51899));
    Odrv4 I__11866 (
            .O(N__51899),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__11865 (
            .O(N__51896),
            .I(N__51890));
    InMux I__11864 (
            .O(N__51895),
            .I(N__51890));
    LocalMux I__11863 (
            .O(N__51890),
            .I(N__51887));
    Odrv12 I__11862 (
            .O(N__51887),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    CascadeMux I__11861 (
            .O(N__51884),
            .I(N__51881));
    InMux I__11860 (
            .O(N__51881),
            .I(N__51878));
    LocalMux I__11859 (
            .O(N__51878),
            .I(N__51874));
    InMux I__11858 (
            .O(N__51877),
            .I(N__51871));
    Span4Mux_v I__11857 (
            .O(N__51874),
            .I(N__51866));
    LocalMux I__11856 (
            .O(N__51871),
            .I(N__51866));
    Odrv4 I__11855 (
            .O(N__51866),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__11854 (
            .O(N__51863),
            .I(N__51860));
    LocalMux I__11853 (
            .O(N__51860),
            .I(N__51856));
    InMux I__11852 (
            .O(N__51859),
            .I(N__51853));
    Span4Mux_v I__11851 (
            .O(N__51856),
            .I(N__51850));
    LocalMux I__11850 (
            .O(N__51853),
            .I(N__51847));
    Odrv4 I__11849 (
            .O(N__51850),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    Odrv4 I__11848 (
            .O(N__51847),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__11847 (
            .O(N__51842),
            .I(N__51836));
    InMux I__11846 (
            .O(N__51841),
            .I(N__51836));
    LocalMux I__11845 (
            .O(N__51836),
            .I(N__51833));
    Odrv4 I__11844 (
            .O(N__51833),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__11843 (
            .O(N__51830),
            .I(N__51824));
    InMux I__11842 (
            .O(N__51829),
            .I(N__51824));
    LocalMux I__11841 (
            .O(N__51824),
            .I(N__51821));
    Odrv12 I__11840 (
            .O(N__51821),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    CascadeMux I__11839 (
            .O(N__51818),
            .I(N__51815));
    InMux I__11838 (
            .O(N__51815),
            .I(N__51810));
    InMux I__11837 (
            .O(N__51814),
            .I(N__51805));
    InMux I__11836 (
            .O(N__51813),
            .I(N__51805));
    LocalMux I__11835 (
            .O(N__51810),
            .I(N__51801));
    LocalMux I__11834 (
            .O(N__51805),
            .I(N__51798));
    InMux I__11833 (
            .O(N__51804),
            .I(N__51795));
    Span4Mux_h I__11832 (
            .O(N__51801),
            .I(N__51790));
    Span4Mux_h I__11831 (
            .O(N__51798),
            .I(N__51790));
    LocalMux I__11830 (
            .O(N__51795),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__11829 (
            .O(N__51790),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__11828 (
            .O(N__51785),
            .I(N__51782));
    InMux I__11827 (
            .O(N__51782),
            .I(N__51777));
    InMux I__11826 (
            .O(N__51781),
            .I(N__51772));
    InMux I__11825 (
            .O(N__51780),
            .I(N__51772));
    LocalMux I__11824 (
            .O(N__51777),
            .I(N__51768));
    LocalMux I__11823 (
            .O(N__51772),
            .I(N__51765));
    InMux I__11822 (
            .O(N__51771),
            .I(N__51762));
    Span4Mux_h I__11821 (
            .O(N__51768),
            .I(N__51757));
    Span4Mux_h I__11820 (
            .O(N__51765),
            .I(N__51757));
    LocalMux I__11819 (
            .O(N__51762),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__11818 (
            .O(N__51757),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    CascadeMux I__11817 (
            .O(N__51752),
            .I(N__51749));
    InMux I__11816 (
            .O(N__51749),
            .I(N__51743));
    InMux I__11815 (
            .O(N__51748),
            .I(N__51740));
    InMux I__11814 (
            .O(N__51747),
            .I(N__51737));
    InMux I__11813 (
            .O(N__51746),
            .I(N__51734));
    LocalMux I__11812 (
            .O(N__51743),
            .I(N__51731));
    LocalMux I__11811 (
            .O(N__51740),
            .I(N__51728));
    LocalMux I__11810 (
            .O(N__51737),
            .I(N__51723));
    LocalMux I__11809 (
            .O(N__51734),
            .I(N__51723));
    Span4Mux_v I__11808 (
            .O(N__51731),
            .I(N__51720));
    Span4Mux_v I__11807 (
            .O(N__51728),
            .I(N__51717));
    Span4Mux_h I__11806 (
            .O(N__51723),
            .I(N__51714));
    Odrv4 I__11805 (
            .O(N__51720),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__11804 (
            .O(N__51717),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__11803 (
            .O(N__51714),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__11802 (
            .O(N__51707),
            .I(N__51702));
    CascadeMux I__11801 (
            .O(N__51706),
            .I(N__51699));
    InMux I__11800 (
            .O(N__51705),
            .I(N__51696));
    InMux I__11799 (
            .O(N__51702),
            .I(N__51693));
    InMux I__11798 (
            .O(N__51699),
            .I(N__51690));
    LocalMux I__11797 (
            .O(N__51696),
            .I(N__51684));
    LocalMux I__11796 (
            .O(N__51693),
            .I(N__51684));
    LocalMux I__11795 (
            .O(N__51690),
            .I(N__51681));
    InMux I__11794 (
            .O(N__51689),
            .I(N__51678));
    Span4Mux_h I__11793 (
            .O(N__51684),
            .I(N__51675));
    Odrv4 I__11792 (
            .O(N__51681),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__11791 (
            .O(N__51678),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__11790 (
            .O(N__51675),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__11789 (
            .O(N__51668),
            .I(N__51665));
    InMux I__11788 (
            .O(N__51665),
            .I(N__51661));
    InMux I__11787 (
            .O(N__51664),
            .I(N__51657));
    LocalMux I__11786 (
            .O(N__51661),
            .I(N__51653));
    InMux I__11785 (
            .O(N__51660),
            .I(N__51650));
    LocalMux I__11784 (
            .O(N__51657),
            .I(N__51647));
    InMux I__11783 (
            .O(N__51656),
            .I(N__51644));
    Span4Mux_h I__11782 (
            .O(N__51653),
            .I(N__51641));
    LocalMux I__11781 (
            .O(N__51650),
            .I(N__51638));
    Odrv12 I__11780 (
            .O(N__51647),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__11779 (
            .O(N__51644),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__11778 (
            .O(N__51641),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__11777 (
            .O(N__51638),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__11776 (
            .O(N__51629),
            .I(N__51623));
    InMux I__11775 (
            .O(N__51628),
            .I(N__51623));
    LocalMux I__11774 (
            .O(N__51623),
            .I(N__51619));
    InMux I__11773 (
            .O(N__51622),
            .I(N__51615));
    Span4Mux_v I__11772 (
            .O(N__51619),
            .I(N__51612));
    InMux I__11771 (
            .O(N__51618),
            .I(N__51609));
    LocalMux I__11770 (
            .O(N__51615),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__11769 (
            .O(N__51612),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__11768 (
            .O(N__51609),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    CascadeMux I__11767 (
            .O(N__51602),
            .I(N__51599));
    InMux I__11766 (
            .O(N__51599),
            .I(N__51596));
    LocalMux I__11765 (
            .O(N__51596),
            .I(N__51590));
    InMux I__11764 (
            .O(N__51595),
            .I(N__51587));
    InMux I__11763 (
            .O(N__51594),
            .I(N__51582));
    InMux I__11762 (
            .O(N__51593),
            .I(N__51582));
    Span4Mux_v I__11761 (
            .O(N__51590),
            .I(N__51579));
    LocalMux I__11760 (
            .O(N__51587),
            .I(N__51576));
    LocalMux I__11759 (
            .O(N__51582),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__11758 (
            .O(N__51579),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__11757 (
            .O(N__51576),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__11756 (
            .O(N__51569),
            .I(N__51566));
    InMux I__11755 (
            .O(N__51566),
            .I(N__51563));
    LocalMux I__11754 (
            .O(N__51563),
            .I(N__51559));
    CascadeMux I__11753 (
            .O(N__51562),
            .I(N__51556));
    Span4Mux_v I__11752 (
            .O(N__51559),
            .I(N__51552));
    InMux I__11751 (
            .O(N__51556),
            .I(N__51549));
    InMux I__11750 (
            .O(N__51555),
            .I(N__51546));
    Odrv4 I__11749 (
            .O(N__51552),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__11748 (
            .O(N__51549),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__11747 (
            .O(N__51546),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__11746 (
            .O(N__51539),
            .I(N__51536));
    LocalMux I__11745 (
            .O(N__51536),
            .I(N__51531));
    CascadeMux I__11744 (
            .O(N__51535),
            .I(N__51528));
    InMux I__11743 (
            .O(N__51534),
            .I(N__51525));
    Span4Mux_h I__11742 (
            .O(N__51531),
            .I(N__51522));
    InMux I__11741 (
            .O(N__51528),
            .I(N__51519));
    LocalMux I__11740 (
            .O(N__51525),
            .I(N__51515));
    Span4Mux_v I__11739 (
            .O(N__51522),
            .I(N__51510));
    LocalMux I__11738 (
            .O(N__51519),
            .I(N__51510));
    InMux I__11737 (
            .O(N__51518),
            .I(N__51507));
    Odrv4 I__11736 (
            .O(N__51515),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__11735 (
            .O(N__51510),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__11734 (
            .O(N__51507),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__11733 (
            .O(N__51500),
            .I(N__51497));
    InMux I__11732 (
            .O(N__51497),
            .I(N__51492));
    InMux I__11731 (
            .O(N__51496),
            .I(N__51489));
    InMux I__11730 (
            .O(N__51495),
            .I(N__51486));
    LocalMux I__11729 (
            .O(N__51492),
            .I(N__51483));
    LocalMux I__11728 (
            .O(N__51489),
            .I(N__51478));
    LocalMux I__11727 (
            .O(N__51486),
            .I(N__51478));
    Span4Mux_h I__11726 (
            .O(N__51483),
            .I(N__51475));
    Span12Mux_s8_v I__11725 (
            .O(N__51478),
            .I(N__51471));
    Span4Mux_h I__11724 (
            .O(N__51475),
            .I(N__51468));
    InMux I__11723 (
            .O(N__51474),
            .I(N__51465));
    Odrv12 I__11722 (
            .O(N__51471),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__11721 (
            .O(N__51468),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__11720 (
            .O(N__51465),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    CascadeMux I__11719 (
            .O(N__51458),
            .I(\current_shift_inst.PI_CTRL.N_77_cascade_ ));
    InMux I__11718 (
            .O(N__51455),
            .I(N__51452));
    LocalMux I__11717 (
            .O(N__51452),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ));
    InMux I__11716 (
            .O(N__51449),
            .I(N__51446));
    LocalMux I__11715 (
            .O(N__51446),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    CascadeMux I__11714 (
            .O(N__51443),
            .I(N__51440));
    InMux I__11713 (
            .O(N__51440),
            .I(N__51437));
    LocalMux I__11712 (
            .O(N__51437),
            .I(N__51433));
    InMux I__11711 (
            .O(N__51436),
            .I(N__51428));
    Span4Mux_h I__11710 (
            .O(N__51433),
            .I(N__51425));
    InMux I__11709 (
            .O(N__51432),
            .I(N__51422));
    InMux I__11708 (
            .O(N__51431),
            .I(N__51419));
    LocalMux I__11707 (
            .O(N__51428),
            .I(N__51416));
    Odrv4 I__11706 (
            .O(N__51425),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__11705 (
            .O(N__51422),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__11704 (
            .O(N__51419),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv12 I__11703 (
            .O(N__51416),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__11702 (
            .O(N__51407),
            .I(N__51404));
    LocalMux I__11701 (
            .O(N__51404),
            .I(\current_shift_inst.PI_CTRL.N_46_16 ));
    InMux I__11700 (
            .O(N__51401),
            .I(N__51398));
    LocalMux I__11699 (
            .O(N__51398),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ));
    InMux I__11698 (
            .O(N__51395),
            .I(N__51392));
    LocalMux I__11697 (
            .O(N__51392),
            .I(N__51389));
    Span4Mux_s3_v I__11696 (
            .O(N__51389),
            .I(N__51386));
    Odrv4 I__11695 (
            .O(N__51386),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    CascadeMux I__11694 (
            .O(N__51383),
            .I(N__51380));
    InMux I__11693 (
            .O(N__51380),
            .I(N__51374));
    InMux I__11692 (
            .O(N__51379),
            .I(N__51371));
    InMux I__11691 (
            .O(N__51378),
            .I(N__51368));
    CascadeMux I__11690 (
            .O(N__51377),
            .I(N__51365));
    LocalMux I__11689 (
            .O(N__51374),
            .I(N__51362));
    LocalMux I__11688 (
            .O(N__51371),
            .I(N__51359));
    LocalMux I__11687 (
            .O(N__51368),
            .I(N__51356));
    InMux I__11686 (
            .O(N__51365),
            .I(N__51353));
    Span4Mux_v I__11685 (
            .O(N__51362),
            .I(N__51346));
    Span4Mux_h I__11684 (
            .O(N__51359),
            .I(N__51346));
    Span4Mux_v I__11683 (
            .O(N__51356),
            .I(N__51346));
    LocalMux I__11682 (
            .O(N__51353),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__11681 (
            .O(N__51346),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__11680 (
            .O(N__51341),
            .I(N__51338));
    LocalMux I__11679 (
            .O(N__51338),
            .I(N__51335));
    Odrv12 I__11678 (
            .O(N__51335),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__11677 (
            .O(N__51332),
            .I(N__51328));
    CascadeMux I__11676 (
            .O(N__51331),
            .I(N__51325));
    InMux I__11675 (
            .O(N__51328),
            .I(N__51321));
    InMux I__11674 (
            .O(N__51325),
            .I(N__51316));
    InMux I__11673 (
            .O(N__51324),
            .I(N__51316));
    LocalMux I__11672 (
            .O(N__51321),
            .I(N__51312));
    LocalMux I__11671 (
            .O(N__51316),
            .I(N__51309));
    InMux I__11670 (
            .O(N__51315),
            .I(N__51306));
    Span4Mux_h I__11669 (
            .O(N__51312),
            .I(N__51301));
    Span4Mux_v I__11668 (
            .O(N__51309),
            .I(N__51301));
    LocalMux I__11667 (
            .O(N__51306),
            .I(N__51298));
    Odrv4 I__11666 (
            .O(N__51301),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__11665 (
            .O(N__51298),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__11664 (
            .O(N__51293),
            .I(N__51290));
    LocalMux I__11663 (
            .O(N__51290),
            .I(N__51287));
    Span4Mux_v I__11662 (
            .O(N__51287),
            .I(N__51284));
    Odrv4 I__11661 (
            .O(N__51284),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    CascadeMux I__11660 (
            .O(N__51281),
            .I(N__51277));
    CascadeMux I__11659 (
            .O(N__51280),
            .I(N__51272));
    InMux I__11658 (
            .O(N__51277),
            .I(N__51269));
    InMux I__11657 (
            .O(N__51276),
            .I(N__51264));
    InMux I__11656 (
            .O(N__51275),
            .I(N__51264));
    InMux I__11655 (
            .O(N__51272),
            .I(N__51261));
    LocalMux I__11654 (
            .O(N__51269),
            .I(N__51254));
    LocalMux I__11653 (
            .O(N__51264),
            .I(N__51254));
    LocalMux I__11652 (
            .O(N__51261),
            .I(N__51254));
    Span4Mux_v I__11651 (
            .O(N__51254),
            .I(N__51251));
    Odrv4 I__11650 (
            .O(N__51251),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__11649 (
            .O(N__51248),
            .I(N__51245));
    LocalMux I__11648 (
            .O(N__51245),
            .I(N__51242));
    Odrv4 I__11647 (
            .O(N__51242),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    CascadeMux I__11646 (
            .O(N__51239),
            .I(N__51236));
    InMux I__11645 (
            .O(N__51236),
            .I(N__51233));
    LocalMux I__11644 (
            .O(N__51233),
            .I(N__51227));
    InMux I__11643 (
            .O(N__51232),
            .I(N__51224));
    InMux I__11642 (
            .O(N__51231),
            .I(N__51219));
    InMux I__11641 (
            .O(N__51230),
            .I(N__51219));
    Odrv4 I__11640 (
            .O(N__51227),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__11639 (
            .O(N__51224),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__11638 (
            .O(N__51219),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__11637 (
            .O(N__51212),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__11636 (
            .O(N__51209),
            .I(N__51206));
    LocalMux I__11635 (
            .O(N__51206),
            .I(N__51203));
    Odrv4 I__11634 (
            .O(N__51203),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ));
    CascadeMux I__11633 (
            .O(N__51200),
            .I(N__51197));
    InMux I__11632 (
            .O(N__51197),
            .I(N__51193));
    CascadeMux I__11631 (
            .O(N__51196),
            .I(N__51190));
    LocalMux I__11630 (
            .O(N__51193),
            .I(N__51185));
    InMux I__11629 (
            .O(N__51190),
            .I(N__51182));
    InMux I__11628 (
            .O(N__51189),
            .I(N__51179));
    InMux I__11627 (
            .O(N__51188),
            .I(N__51176));
    Odrv4 I__11626 (
            .O(N__51185),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__11625 (
            .O(N__51182),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__11624 (
            .O(N__51179),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__11623 (
            .O(N__51176),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__11622 (
            .O(N__51167),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__11621 (
            .O(N__51164),
            .I(N__51161));
    LocalMux I__11620 (
            .O(N__51161),
            .I(N__51158));
    Span4Mux_v I__11619 (
            .O(N__51158),
            .I(N__51155));
    Odrv4 I__11618 (
            .O(N__51155),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ));
    CascadeMux I__11617 (
            .O(N__51152),
            .I(N__51149));
    InMux I__11616 (
            .O(N__51149),
            .I(N__51145));
    CascadeMux I__11615 (
            .O(N__51148),
            .I(N__51142));
    LocalMux I__11614 (
            .O(N__51145),
            .I(N__51137));
    InMux I__11613 (
            .O(N__51142),
            .I(N__51134));
    InMux I__11612 (
            .O(N__51141),
            .I(N__51131));
    InMux I__11611 (
            .O(N__51140),
            .I(N__51128));
    Odrv12 I__11610 (
            .O(N__51137),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__11609 (
            .O(N__51134),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__11608 (
            .O(N__51131),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__11607 (
            .O(N__51128),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__11606 (
            .O(N__51119),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__11605 (
            .O(N__51116),
            .I(N__51113));
    LocalMux I__11604 (
            .O(N__51113),
            .I(N__51110));
    Span4Mux_h I__11603 (
            .O(N__51110),
            .I(N__51107));
    Odrv4 I__11602 (
            .O(N__51107),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ));
    CascadeMux I__11601 (
            .O(N__51104),
            .I(N__51101));
    InMux I__11600 (
            .O(N__51101),
            .I(N__51097));
    CascadeMux I__11599 (
            .O(N__51100),
            .I(N__51093));
    LocalMux I__11598 (
            .O(N__51097),
            .I(N__51089));
    InMux I__11597 (
            .O(N__51096),
            .I(N__51086));
    InMux I__11596 (
            .O(N__51093),
            .I(N__51081));
    InMux I__11595 (
            .O(N__51092),
            .I(N__51081));
    Odrv12 I__11594 (
            .O(N__51089),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__11593 (
            .O(N__51086),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__11592 (
            .O(N__51081),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__11591 (
            .O(N__51074),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__11590 (
            .O(N__51071),
            .I(N__51067));
    CascadeMux I__11589 (
            .O(N__51070),
            .I(N__51064));
    LocalMux I__11588 (
            .O(N__51067),
            .I(N__51059));
    InMux I__11587 (
            .O(N__51064),
            .I(N__51056));
    InMux I__11586 (
            .O(N__51063),
            .I(N__51053));
    InMux I__11585 (
            .O(N__51062),
            .I(N__51050));
    Odrv12 I__11584 (
            .O(N__51059),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__11583 (
            .O(N__51056),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__11582 (
            .O(N__51053),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__11581 (
            .O(N__51050),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__11580 (
            .O(N__51041),
            .I(N__51038));
    InMux I__11579 (
            .O(N__51038),
            .I(N__51035));
    LocalMux I__11578 (
            .O(N__51035),
            .I(N__51032));
    Span4Mux_v I__11577 (
            .O(N__51032),
            .I(N__51029));
    Odrv4 I__11576 (
            .O(N__51029),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ));
    InMux I__11575 (
            .O(N__51026),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__11574 (
            .O(N__51023),
            .I(N__51020));
    LocalMux I__11573 (
            .O(N__51020),
            .I(N__51017));
    Odrv4 I__11572 (
            .O(N__51017),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ));
    InMux I__11571 (
            .O(N__51014),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    CascadeMux I__11570 (
            .O(N__51011),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__11569 (
            .O(N__51008),
            .I(N__51005));
    LocalMux I__11568 (
            .O(N__51005),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    InMux I__11567 (
            .O(N__51002),
            .I(N__50999));
    LocalMux I__11566 (
            .O(N__50999),
            .I(N__50996));
    Odrv4 I__11565 (
            .O(N__50996),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    InMux I__11564 (
            .O(N__50993),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__11563 (
            .O(N__50990),
            .I(N__50987));
    LocalMux I__11562 (
            .O(N__50987),
            .I(N__50984));
    Span12Mux_s7_v I__11561 (
            .O(N__50984),
            .I(N__50981));
    Odrv12 I__11560 (
            .O(N__50981),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    InMux I__11559 (
            .O(N__50978),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__11558 (
            .O(N__50975),
            .I(N__50972));
    LocalMux I__11557 (
            .O(N__50972),
            .I(N__50969));
    Odrv4 I__11556 (
            .O(N__50969),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    InMux I__11555 (
            .O(N__50966),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__11554 (
            .O(N__50963),
            .I(N__50960));
    LocalMux I__11553 (
            .O(N__50960),
            .I(N__50957));
    Odrv4 I__11552 (
            .O(N__50957),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    CascadeMux I__11551 (
            .O(N__50954),
            .I(N__50951));
    InMux I__11550 (
            .O(N__50951),
            .I(N__50946));
    InMux I__11549 (
            .O(N__50950),
            .I(N__50940));
    InMux I__11548 (
            .O(N__50949),
            .I(N__50940));
    LocalMux I__11547 (
            .O(N__50946),
            .I(N__50937));
    InMux I__11546 (
            .O(N__50945),
            .I(N__50934));
    LocalMux I__11545 (
            .O(N__50940),
            .I(N__50931));
    Odrv4 I__11544 (
            .O(N__50937),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__11543 (
            .O(N__50934),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__11542 (
            .O(N__50931),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__11541 (
            .O(N__50924),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    CascadeMux I__11540 (
            .O(N__50921),
            .I(N__50918));
    InMux I__11539 (
            .O(N__50918),
            .I(N__50915));
    LocalMux I__11538 (
            .O(N__50915),
            .I(N__50912));
    Odrv4 I__11537 (
            .O(N__50912),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    InMux I__11536 (
            .O(N__50909),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__11535 (
            .O(N__50906),
            .I(N__50900));
    InMux I__11534 (
            .O(N__50905),
            .I(N__50897));
    InMux I__11533 (
            .O(N__50904),
            .I(N__50892));
    InMux I__11532 (
            .O(N__50903),
            .I(N__50892));
    LocalMux I__11531 (
            .O(N__50900),
            .I(N__50889));
    LocalMux I__11530 (
            .O(N__50897),
            .I(N__50884));
    LocalMux I__11529 (
            .O(N__50892),
            .I(N__50884));
    Odrv4 I__11528 (
            .O(N__50889),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__11527 (
            .O(N__50884),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__11526 (
            .O(N__50879),
            .I(N__50876));
    InMux I__11525 (
            .O(N__50876),
            .I(N__50873));
    LocalMux I__11524 (
            .O(N__50873),
            .I(N__50870));
    Span4Mux_h I__11523 (
            .O(N__50870),
            .I(N__50867));
    Odrv4 I__11522 (
            .O(N__50867),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    InMux I__11521 (
            .O(N__50864),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__11520 (
            .O(N__50861),
            .I(N__50858));
    LocalMux I__11519 (
            .O(N__50858),
            .I(N__50855));
    Span4Mux_h I__11518 (
            .O(N__50855),
            .I(N__50852));
    Odrv4 I__11517 (
            .O(N__50852),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    CascadeMux I__11516 (
            .O(N__50849),
            .I(N__50845));
    CascadeMux I__11515 (
            .O(N__50848),
            .I(N__50841));
    InMux I__11514 (
            .O(N__50845),
            .I(N__50837));
    CascadeMux I__11513 (
            .O(N__50844),
            .I(N__50834));
    InMux I__11512 (
            .O(N__50841),
            .I(N__50829));
    InMux I__11511 (
            .O(N__50840),
            .I(N__50829));
    LocalMux I__11510 (
            .O(N__50837),
            .I(N__50826));
    InMux I__11509 (
            .O(N__50834),
            .I(N__50823));
    LocalMux I__11508 (
            .O(N__50829),
            .I(N__50820));
    Odrv12 I__11507 (
            .O(N__50826),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__11506 (
            .O(N__50823),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__11505 (
            .O(N__50820),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__11504 (
            .O(N__50813),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    InMux I__11503 (
            .O(N__50810),
            .I(N__50807));
    LocalMux I__11502 (
            .O(N__50807),
            .I(N__50804));
    Odrv4 I__11501 (
            .O(N__50804),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    CascadeMux I__11500 (
            .O(N__50801),
            .I(N__50798));
    InMux I__11499 (
            .O(N__50798),
            .I(N__50795));
    LocalMux I__11498 (
            .O(N__50795),
            .I(N__50790));
    CascadeMux I__11497 (
            .O(N__50794),
            .I(N__50787));
    CascadeMux I__11496 (
            .O(N__50793),
            .I(N__50783));
    Span4Mux_h I__11495 (
            .O(N__50790),
            .I(N__50780));
    InMux I__11494 (
            .O(N__50787),
            .I(N__50777));
    InMux I__11493 (
            .O(N__50786),
            .I(N__50772));
    InMux I__11492 (
            .O(N__50783),
            .I(N__50772));
    Odrv4 I__11491 (
            .O(N__50780),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__11490 (
            .O(N__50777),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__11489 (
            .O(N__50772),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__11488 (
            .O(N__50765),
            .I(bfn_18_26_0_));
    InMux I__11487 (
            .O(N__50762),
            .I(N__50759));
    LocalMux I__11486 (
            .O(N__50759),
            .I(N__50756));
    Odrv4 I__11485 (
            .O(N__50756),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__11484 (
            .O(N__50753),
            .I(N__50750));
    InMux I__11483 (
            .O(N__50750),
            .I(N__50744));
    InMux I__11482 (
            .O(N__50749),
            .I(N__50741));
    InMux I__11481 (
            .O(N__50748),
            .I(N__50736));
    InMux I__11480 (
            .O(N__50747),
            .I(N__50736));
    LocalMux I__11479 (
            .O(N__50744),
            .I(N__50731));
    LocalMux I__11478 (
            .O(N__50741),
            .I(N__50731));
    LocalMux I__11477 (
            .O(N__50736),
            .I(N__50728));
    Span4Mux_h I__11476 (
            .O(N__50731),
            .I(N__50725));
    Odrv4 I__11475 (
            .O(N__50728),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__11474 (
            .O(N__50725),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__11473 (
            .O(N__50720),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__11472 (
            .O(N__50717),
            .I(N__50714));
    LocalMux I__11471 (
            .O(N__50714),
            .I(N__50711));
    Odrv12 I__11470 (
            .O(N__50711),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__11469 (
            .O(N__50708),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__11468 (
            .O(N__50705),
            .I(N__50702));
    LocalMux I__11467 (
            .O(N__50702),
            .I(N__50699));
    Odrv12 I__11466 (
            .O(N__50699),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    CascadeMux I__11465 (
            .O(N__50696),
            .I(N__50693));
    InMux I__11464 (
            .O(N__50693),
            .I(N__50689));
    CascadeMux I__11463 (
            .O(N__50692),
            .I(N__50686));
    LocalMux I__11462 (
            .O(N__50689),
            .I(N__50682));
    InMux I__11461 (
            .O(N__50686),
            .I(N__50678));
    InMux I__11460 (
            .O(N__50685),
            .I(N__50675));
    Span4Mux_h I__11459 (
            .O(N__50682),
            .I(N__50672));
    CascadeMux I__11458 (
            .O(N__50681),
            .I(N__50669));
    LocalMux I__11457 (
            .O(N__50678),
            .I(N__50664));
    LocalMux I__11456 (
            .O(N__50675),
            .I(N__50664));
    Span4Mux_v I__11455 (
            .O(N__50672),
            .I(N__50661));
    InMux I__11454 (
            .O(N__50669),
            .I(N__50658));
    Span12Mux_v I__11453 (
            .O(N__50664),
            .I(N__50655));
    Odrv4 I__11452 (
            .O(N__50661),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__11451 (
            .O(N__50658),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv12 I__11450 (
            .O(N__50655),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__11449 (
            .O(N__50648),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__11448 (
            .O(N__50645),
            .I(N__50642));
    LocalMux I__11447 (
            .O(N__50642),
            .I(N__50639));
    Odrv12 I__11446 (
            .O(N__50639),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__11445 (
            .O(N__50636),
            .I(N__50633));
    InMux I__11444 (
            .O(N__50633),
            .I(N__50630));
    LocalMux I__11443 (
            .O(N__50630),
            .I(N__50626));
    InMux I__11442 (
            .O(N__50629),
            .I(N__50623));
    Span4Mux_h I__11441 (
            .O(N__50626),
            .I(N__50619));
    LocalMux I__11440 (
            .O(N__50623),
            .I(N__50615));
    InMux I__11439 (
            .O(N__50622),
            .I(N__50612));
    Span4Mux_v I__11438 (
            .O(N__50619),
            .I(N__50609));
    InMux I__11437 (
            .O(N__50618),
            .I(N__50606));
    Span4Mux_v I__11436 (
            .O(N__50615),
            .I(N__50603));
    LocalMux I__11435 (
            .O(N__50612),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__11434 (
            .O(N__50609),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__11433 (
            .O(N__50606),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__11432 (
            .O(N__50603),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__11431 (
            .O(N__50594),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__11430 (
            .O(N__50591),
            .I(N__50588));
    LocalMux I__11429 (
            .O(N__50588),
            .I(N__50585));
    Odrv4 I__11428 (
            .O(N__50585),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__11427 (
            .O(N__50582),
            .I(N__50579));
    InMux I__11426 (
            .O(N__50579),
            .I(N__50575));
    InMux I__11425 (
            .O(N__50578),
            .I(N__50572));
    LocalMux I__11424 (
            .O(N__50575),
            .I(N__50565));
    LocalMux I__11423 (
            .O(N__50572),
            .I(N__50565));
    InMux I__11422 (
            .O(N__50571),
            .I(N__50562));
    InMux I__11421 (
            .O(N__50570),
            .I(N__50559));
    Span4Mux_h I__11420 (
            .O(N__50565),
            .I(N__50556));
    LocalMux I__11419 (
            .O(N__50562),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__11418 (
            .O(N__50559),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__11417 (
            .O(N__50556),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__11416 (
            .O(N__50549),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__11415 (
            .O(N__50546),
            .I(N__50543));
    LocalMux I__11414 (
            .O(N__50543),
            .I(N__50540));
    Span4Mux_h I__11413 (
            .O(N__50540),
            .I(N__50537));
    Odrv4 I__11412 (
            .O(N__50537),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__11411 (
            .O(N__50534),
            .I(N__50531));
    InMux I__11410 (
            .O(N__50531),
            .I(N__50528));
    LocalMux I__11409 (
            .O(N__50528),
            .I(N__50523));
    InMux I__11408 (
            .O(N__50527),
            .I(N__50517));
    InMux I__11407 (
            .O(N__50526),
            .I(N__50517));
    Span4Mux_v I__11406 (
            .O(N__50523),
            .I(N__50514));
    InMux I__11405 (
            .O(N__50522),
            .I(N__50511));
    LocalMux I__11404 (
            .O(N__50517),
            .I(N__50508));
    Odrv4 I__11403 (
            .O(N__50514),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__11402 (
            .O(N__50511),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__11401 (
            .O(N__50508),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__11400 (
            .O(N__50501),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__11399 (
            .O(N__50498),
            .I(N__50495));
    LocalMux I__11398 (
            .O(N__50495),
            .I(N__50492));
    Odrv12 I__11397 (
            .O(N__50492),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__11396 (
            .O(N__50489),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    InMux I__11395 (
            .O(N__50486),
            .I(N__50483));
    LocalMux I__11394 (
            .O(N__50483),
            .I(N__50480));
    Span4Mux_h I__11393 (
            .O(N__50480),
            .I(N__50477));
    Span4Mux_h I__11392 (
            .O(N__50477),
            .I(N__50474));
    Odrv4 I__11391 (
            .O(N__50474),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    InMux I__11390 (
            .O(N__50471),
            .I(bfn_18_25_0_));
    InMux I__11389 (
            .O(N__50468),
            .I(N__50465));
    LocalMux I__11388 (
            .O(N__50465),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__11387 (
            .O(N__50462),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    CascadeMux I__11386 (
            .O(N__50459),
            .I(N__50456));
    InMux I__11385 (
            .O(N__50456),
            .I(N__50453));
    LocalMux I__11384 (
            .O(N__50453),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__11383 (
            .O(N__50450),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__11382 (
            .O(N__50447),
            .I(N__50444));
    LocalMux I__11381 (
            .O(N__50444),
            .I(N__50441));
    Odrv4 I__11380 (
            .O(N__50441),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__11379 (
            .O(N__50438),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__11378 (
            .O(N__50435),
            .I(N__50432));
    LocalMux I__11377 (
            .O(N__50432),
            .I(N__50429));
    Span4Mux_h I__11376 (
            .O(N__50429),
            .I(N__50426));
    Odrv4 I__11375 (
            .O(N__50426),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__11374 (
            .O(N__50423),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__11373 (
            .O(N__50420),
            .I(N__50417));
    LocalMux I__11372 (
            .O(N__50417),
            .I(N__50414));
    Odrv12 I__11371 (
            .O(N__50414),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__11370 (
            .O(N__50411),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__11369 (
            .O(N__50408),
            .I(N__50405));
    LocalMux I__11368 (
            .O(N__50405),
            .I(N__50402));
    Odrv12 I__11367 (
            .O(N__50402),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__11366 (
            .O(N__50399),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__11365 (
            .O(N__50396),
            .I(N__50393));
    LocalMux I__11364 (
            .O(N__50393),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__11363 (
            .O(N__50390),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    InMux I__11362 (
            .O(N__50387),
            .I(N__50384));
    LocalMux I__11361 (
            .O(N__50384),
            .I(N__50381));
    Odrv4 I__11360 (
            .O(N__50381),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__11359 (
            .O(N__50378),
            .I(bfn_18_24_0_));
    InMux I__11358 (
            .O(N__50375),
            .I(N__50371));
    InMux I__11357 (
            .O(N__50374),
            .I(N__50368));
    LocalMux I__11356 (
            .O(N__50371),
            .I(N__50365));
    LocalMux I__11355 (
            .O(N__50368),
            .I(N__50360));
    Span12Mux_s8_v I__11354 (
            .O(N__50365),
            .I(N__50360));
    Odrv12 I__11353 (
            .O(N__50360),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__11352 (
            .O(N__50357),
            .I(N__50354));
    LocalMux I__11351 (
            .O(N__50354),
            .I(N__50350));
    InMux I__11350 (
            .O(N__50353),
            .I(N__50347));
    Span4Mux_v I__11349 (
            .O(N__50350),
            .I(N__50344));
    LocalMux I__11348 (
            .O(N__50347),
            .I(N__50339));
    Span4Mux_h I__11347 (
            .O(N__50344),
            .I(N__50339));
    Span4Mux_h I__11346 (
            .O(N__50339),
            .I(N__50336));
    Odrv4 I__11345 (
            .O(N__50336),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__11344 (
            .O(N__50333),
            .I(N__50330));
    LocalMux I__11343 (
            .O(N__50330),
            .I(N__50326));
    InMux I__11342 (
            .O(N__50329),
            .I(N__50323));
    Span4Mux_s2_h I__11341 (
            .O(N__50326),
            .I(N__50320));
    LocalMux I__11340 (
            .O(N__50323),
            .I(N__50315));
    Span4Mux_h I__11339 (
            .O(N__50320),
            .I(N__50315));
    Span4Mux_v I__11338 (
            .O(N__50315),
            .I(N__50312));
    Odrv4 I__11337 (
            .O(N__50312),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__11336 (
            .O(N__50309),
            .I(N__50306));
    LocalMux I__11335 (
            .O(N__50306),
            .I(N__50303));
    Span4Mux_s1_h I__11334 (
            .O(N__50303),
            .I(N__50299));
    InMux I__11333 (
            .O(N__50302),
            .I(N__50296));
    Span4Mux_h I__11332 (
            .O(N__50299),
            .I(N__50293));
    LocalMux I__11331 (
            .O(N__50296),
            .I(N__50290));
    Span4Mux_h I__11330 (
            .O(N__50293),
            .I(N__50287));
    Odrv4 I__11329 (
            .O(N__50290),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__11328 (
            .O(N__50287),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__11327 (
            .O(N__50282),
            .I(N__50279));
    LocalMux I__11326 (
            .O(N__50279),
            .I(N__50275));
    InMux I__11325 (
            .O(N__50278),
            .I(N__50272));
    Span4Mux_v I__11324 (
            .O(N__50275),
            .I(N__50269));
    LocalMux I__11323 (
            .O(N__50272),
            .I(N__50264));
    Span4Mux_h I__11322 (
            .O(N__50269),
            .I(N__50264));
    Span4Mux_h I__11321 (
            .O(N__50264),
            .I(N__50261));
    Odrv4 I__11320 (
            .O(N__50261),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__11319 (
            .O(N__50258),
            .I(N__50254));
    InMux I__11318 (
            .O(N__50257),
            .I(N__50251));
    LocalMux I__11317 (
            .O(N__50254),
            .I(N__50248));
    LocalMux I__11316 (
            .O(N__50251),
            .I(N__50245));
    Span12Mux_s10_h I__11315 (
            .O(N__50248),
            .I(N__50242));
    Odrv4 I__11314 (
            .O(N__50245),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv12 I__11313 (
            .O(N__50242),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__11312 (
            .O(N__50237),
            .I(N__50234));
    LocalMux I__11311 (
            .O(N__50234),
            .I(N__50230));
    InMux I__11310 (
            .O(N__50233),
            .I(N__50227));
    Span4Mux_s2_h I__11309 (
            .O(N__50230),
            .I(N__50224));
    LocalMux I__11308 (
            .O(N__50227),
            .I(N__50219));
    Span4Mux_h I__11307 (
            .O(N__50224),
            .I(N__50219));
    Span4Mux_v I__11306 (
            .O(N__50219),
            .I(N__50216));
    Odrv4 I__11305 (
            .O(N__50216),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__11304 (
            .O(N__50213),
            .I(N__50210));
    LocalMux I__11303 (
            .O(N__50210),
            .I(N__50207));
    Span4Mux_s2_h I__11302 (
            .O(N__50207),
            .I(N__50203));
    InMux I__11301 (
            .O(N__50206),
            .I(N__50200));
    Span4Mux_h I__11300 (
            .O(N__50203),
            .I(N__50197));
    LocalMux I__11299 (
            .O(N__50200),
            .I(N__50194));
    Span4Mux_h I__11298 (
            .O(N__50197),
            .I(N__50191));
    Odrv4 I__11297 (
            .O(N__50194),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__11296 (
            .O(N__50191),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__11295 (
            .O(N__50186),
            .I(N__50182));
    InMux I__11294 (
            .O(N__50185),
            .I(N__50179));
    LocalMux I__11293 (
            .O(N__50182),
            .I(N__50176));
    LocalMux I__11292 (
            .O(N__50179),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    Odrv4 I__11291 (
            .O(N__50176),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__11290 (
            .O(N__50171),
            .I(N__50168));
    LocalMux I__11289 (
            .O(N__50168),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ));
    InMux I__11288 (
            .O(N__50165),
            .I(N__50159));
    InMux I__11287 (
            .O(N__50164),
            .I(N__50159));
    LocalMux I__11286 (
            .O(N__50159),
            .I(N__50155));
    InMux I__11285 (
            .O(N__50158),
            .I(N__50152));
    Span4Mux_v I__11284 (
            .O(N__50155),
            .I(N__50149));
    LocalMux I__11283 (
            .O(N__50152),
            .I(N__50146));
    Odrv4 I__11282 (
            .O(N__50149),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__11281 (
            .O(N__50146),
            .I(\current_shift_inst.un4_control_input1_4 ));
    CascadeMux I__11280 (
            .O(N__50141),
            .I(N__50138));
    InMux I__11279 (
            .O(N__50138),
            .I(N__50132));
    InMux I__11278 (
            .O(N__50137),
            .I(N__50127));
    InMux I__11277 (
            .O(N__50136),
            .I(N__50127));
    CascadeMux I__11276 (
            .O(N__50135),
            .I(N__50122));
    LocalMux I__11275 (
            .O(N__50132),
            .I(N__50112));
    LocalMux I__11274 (
            .O(N__50127),
            .I(N__50112));
    CascadeMux I__11273 (
            .O(N__50126),
            .I(N__50108));
    InMux I__11272 (
            .O(N__50125),
            .I(N__50092));
    InMux I__11271 (
            .O(N__50122),
            .I(N__50068));
    InMux I__11270 (
            .O(N__50121),
            .I(N__50068));
    InMux I__11269 (
            .O(N__50120),
            .I(N__50068));
    InMux I__11268 (
            .O(N__50119),
            .I(N__50068));
    InMux I__11267 (
            .O(N__50118),
            .I(N__50068));
    InMux I__11266 (
            .O(N__50117),
            .I(N__50068));
    Span4Mux_h I__11265 (
            .O(N__50112),
            .I(N__50065));
    InMux I__11264 (
            .O(N__50111),
            .I(N__50060));
    InMux I__11263 (
            .O(N__50108),
            .I(N__50060));
    InMux I__11262 (
            .O(N__50107),
            .I(N__50050));
    InMux I__11261 (
            .O(N__50106),
            .I(N__50050));
    InMux I__11260 (
            .O(N__50105),
            .I(N__50050));
    InMux I__11259 (
            .O(N__50104),
            .I(N__50050));
    InMux I__11258 (
            .O(N__50103),
            .I(N__50046));
    InMux I__11257 (
            .O(N__50102),
            .I(N__50033));
    InMux I__11256 (
            .O(N__50101),
            .I(N__50033));
    InMux I__11255 (
            .O(N__50100),
            .I(N__50033));
    InMux I__11254 (
            .O(N__50099),
            .I(N__50033));
    InMux I__11253 (
            .O(N__50098),
            .I(N__50033));
    InMux I__11252 (
            .O(N__50097),
            .I(N__50033));
    InMux I__11251 (
            .O(N__50096),
            .I(N__50028));
    InMux I__11250 (
            .O(N__50095),
            .I(N__50028));
    LocalMux I__11249 (
            .O(N__50092),
            .I(N__50025));
    InMux I__11248 (
            .O(N__50091),
            .I(N__50022));
    InMux I__11247 (
            .O(N__50090),
            .I(N__50004));
    InMux I__11246 (
            .O(N__50089),
            .I(N__50004));
    InMux I__11245 (
            .O(N__50088),
            .I(N__50004));
    InMux I__11244 (
            .O(N__50087),
            .I(N__50004));
    InMux I__11243 (
            .O(N__50086),
            .I(N__50004));
    InMux I__11242 (
            .O(N__50085),
            .I(N__50004));
    InMux I__11241 (
            .O(N__50084),
            .I(N__50004));
    InMux I__11240 (
            .O(N__50083),
            .I(N__50004));
    InMux I__11239 (
            .O(N__50082),
            .I(N__49999));
    InMux I__11238 (
            .O(N__50081),
            .I(N__49999));
    LocalMux I__11237 (
            .O(N__50068),
            .I(N__49982));
    Span4Mux_v I__11236 (
            .O(N__50065),
            .I(N__49973));
    LocalMux I__11235 (
            .O(N__50060),
            .I(N__49973));
    InMux I__11234 (
            .O(N__50059),
            .I(N__49970));
    LocalMux I__11233 (
            .O(N__50050),
            .I(N__49967));
    InMux I__11232 (
            .O(N__50049),
            .I(N__49964));
    LocalMux I__11231 (
            .O(N__50046),
            .I(N__49959));
    LocalMux I__11230 (
            .O(N__50033),
            .I(N__49959));
    LocalMux I__11229 (
            .O(N__50028),
            .I(N__49952));
    Span4Mux_h I__11228 (
            .O(N__50025),
            .I(N__49952));
    LocalMux I__11227 (
            .O(N__50022),
            .I(N__49952));
    CascadeMux I__11226 (
            .O(N__50021),
            .I(N__49937));
    LocalMux I__11225 (
            .O(N__50004),
            .I(N__49930));
    LocalMux I__11224 (
            .O(N__49999),
            .I(N__49930));
    InMux I__11223 (
            .O(N__49998),
            .I(N__49923));
    InMux I__11222 (
            .O(N__49997),
            .I(N__49923));
    InMux I__11221 (
            .O(N__49996),
            .I(N__49923));
    InMux I__11220 (
            .O(N__49995),
            .I(N__49912));
    InMux I__11219 (
            .O(N__49994),
            .I(N__49912));
    InMux I__11218 (
            .O(N__49993),
            .I(N__49912));
    InMux I__11217 (
            .O(N__49992),
            .I(N__49912));
    InMux I__11216 (
            .O(N__49991),
            .I(N__49912));
    InMux I__11215 (
            .O(N__49990),
            .I(N__49899));
    InMux I__11214 (
            .O(N__49989),
            .I(N__49899));
    InMux I__11213 (
            .O(N__49988),
            .I(N__49899));
    InMux I__11212 (
            .O(N__49987),
            .I(N__49899));
    InMux I__11211 (
            .O(N__49986),
            .I(N__49899));
    InMux I__11210 (
            .O(N__49985),
            .I(N__49899));
    Span4Mux_h I__11209 (
            .O(N__49982),
            .I(N__49896));
    InMux I__11208 (
            .O(N__49981),
            .I(N__49887));
    InMux I__11207 (
            .O(N__49980),
            .I(N__49887));
    InMux I__11206 (
            .O(N__49979),
            .I(N__49887));
    InMux I__11205 (
            .O(N__49978),
            .I(N__49887));
    Span4Mux_h I__11204 (
            .O(N__49973),
            .I(N__49884));
    LocalMux I__11203 (
            .O(N__49970),
            .I(N__49881));
    Span4Mux_v I__11202 (
            .O(N__49967),
            .I(N__49878));
    LocalMux I__11201 (
            .O(N__49964),
            .I(N__49871));
    Span4Mux_h I__11200 (
            .O(N__49959),
            .I(N__49871));
    Span4Mux_v I__11199 (
            .O(N__49952),
            .I(N__49871));
    InMux I__11198 (
            .O(N__49951),
            .I(N__49854));
    InMux I__11197 (
            .O(N__49950),
            .I(N__49854));
    InMux I__11196 (
            .O(N__49949),
            .I(N__49854));
    InMux I__11195 (
            .O(N__49948),
            .I(N__49854));
    InMux I__11194 (
            .O(N__49947),
            .I(N__49854));
    InMux I__11193 (
            .O(N__49946),
            .I(N__49854));
    InMux I__11192 (
            .O(N__49945),
            .I(N__49854));
    InMux I__11191 (
            .O(N__49944),
            .I(N__49854));
    InMux I__11190 (
            .O(N__49943),
            .I(N__49851));
    InMux I__11189 (
            .O(N__49942),
            .I(N__49838));
    InMux I__11188 (
            .O(N__49941),
            .I(N__49838));
    InMux I__11187 (
            .O(N__49940),
            .I(N__49838));
    InMux I__11186 (
            .O(N__49937),
            .I(N__49838));
    InMux I__11185 (
            .O(N__49936),
            .I(N__49838));
    InMux I__11184 (
            .O(N__49935),
            .I(N__49838));
    Span12Mux_h I__11183 (
            .O(N__49930),
            .I(N__49835));
    LocalMux I__11182 (
            .O(N__49923),
            .I(N__49824));
    LocalMux I__11181 (
            .O(N__49912),
            .I(N__49824));
    LocalMux I__11180 (
            .O(N__49899),
            .I(N__49824));
    Sp12to4 I__11179 (
            .O(N__49896),
            .I(N__49824));
    LocalMux I__11178 (
            .O(N__49887),
            .I(N__49824));
    Odrv4 I__11177 (
            .O(N__49884),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11176 (
            .O(N__49881),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11175 (
            .O(N__49878),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11174 (
            .O(N__49871),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11173 (
            .O(N__49854),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11172 (
            .O(N__49851),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11171 (
            .O(N__49838),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__11170 (
            .O(N__49835),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__11169 (
            .O(N__49824),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__11168 (
            .O(N__49805),
            .I(N__49801));
    InMux I__11167 (
            .O(N__49804),
            .I(N__49796));
    InMux I__11166 (
            .O(N__49801),
            .I(N__49796));
    LocalMux I__11165 (
            .O(N__49796),
            .I(N__49793));
    Span4Mux_v I__11164 (
            .O(N__49793),
            .I(N__49789));
    InMux I__11163 (
            .O(N__49792),
            .I(N__49786));
    Span4Mux_h I__11162 (
            .O(N__49789),
            .I(N__49782));
    LocalMux I__11161 (
            .O(N__49786),
            .I(N__49779));
    InMux I__11160 (
            .O(N__49785),
            .I(N__49776));
    Odrv4 I__11159 (
            .O(N__49782),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv12 I__11158 (
            .O(N__49779),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__11157 (
            .O(N__49776),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    CascadeMux I__11156 (
            .O(N__49769),
            .I(N__49762));
    CascadeMux I__11155 (
            .O(N__49768),
            .I(N__49753));
    CascadeMux I__11154 (
            .O(N__49767),
            .I(N__49747));
    CascadeMux I__11153 (
            .O(N__49766),
            .I(N__49743));
    CascadeMux I__11152 (
            .O(N__49765),
            .I(N__49740));
    InMux I__11151 (
            .O(N__49762),
            .I(N__49737));
    CascadeMux I__11150 (
            .O(N__49761),
            .I(N__49733));
    CascadeMux I__11149 (
            .O(N__49760),
            .I(N__49730));
    CascadeMux I__11148 (
            .O(N__49759),
            .I(N__49724));
    CascadeMux I__11147 (
            .O(N__49758),
            .I(N__49720));
    CascadeMux I__11146 (
            .O(N__49757),
            .I(N__49709));
    CascadeMux I__11145 (
            .O(N__49756),
            .I(N__49702));
    InMux I__11144 (
            .O(N__49753),
            .I(N__49685));
    InMux I__11143 (
            .O(N__49752),
            .I(N__49685));
    InMux I__11142 (
            .O(N__49751),
            .I(N__49685));
    InMux I__11141 (
            .O(N__49750),
            .I(N__49685));
    InMux I__11140 (
            .O(N__49747),
            .I(N__49685));
    InMux I__11139 (
            .O(N__49746),
            .I(N__49685));
    InMux I__11138 (
            .O(N__49743),
            .I(N__49685));
    InMux I__11137 (
            .O(N__49740),
            .I(N__49685));
    LocalMux I__11136 (
            .O(N__49737),
            .I(N__49682));
    InMux I__11135 (
            .O(N__49736),
            .I(N__49667));
    InMux I__11134 (
            .O(N__49733),
            .I(N__49667));
    InMux I__11133 (
            .O(N__49730),
            .I(N__49667));
    InMux I__11132 (
            .O(N__49729),
            .I(N__49667));
    InMux I__11131 (
            .O(N__49728),
            .I(N__49667));
    InMux I__11130 (
            .O(N__49727),
            .I(N__49667));
    InMux I__11129 (
            .O(N__49724),
            .I(N__49667));
    InMux I__11128 (
            .O(N__49723),
            .I(N__49662));
    InMux I__11127 (
            .O(N__49720),
            .I(N__49662));
    InMux I__11126 (
            .O(N__49719),
            .I(N__49651));
    InMux I__11125 (
            .O(N__49718),
            .I(N__49651));
    InMux I__11124 (
            .O(N__49717),
            .I(N__49651));
    InMux I__11123 (
            .O(N__49716),
            .I(N__49651));
    InMux I__11122 (
            .O(N__49715),
            .I(N__49651));
    InMux I__11121 (
            .O(N__49714),
            .I(N__49640));
    InMux I__11120 (
            .O(N__49713),
            .I(N__49640));
    InMux I__11119 (
            .O(N__49712),
            .I(N__49640));
    InMux I__11118 (
            .O(N__49709),
            .I(N__49640));
    CascadeMux I__11117 (
            .O(N__49708),
            .I(N__49636));
    CascadeMux I__11116 (
            .O(N__49707),
            .I(N__49631));
    CascadeMux I__11115 (
            .O(N__49706),
            .I(N__49628));
    CascadeMux I__11114 (
            .O(N__49705),
            .I(N__49625));
    InMux I__11113 (
            .O(N__49702),
            .I(N__49609));
    LocalMux I__11112 (
            .O(N__49685),
            .I(N__49606));
    Span4Mux_v I__11111 (
            .O(N__49682),
            .I(N__49597));
    LocalMux I__11110 (
            .O(N__49667),
            .I(N__49597));
    LocalMux I__11109 (
            .O(N__49662),
            .I(N__49597));
    LocalMux I__11108 (
            .O(N__49651),
            .I(N__49597));
    InMux I__11107 (
            .O(N__49650),
            .I(N__49592));
    InMux I__11106 (
            .O(N__49649),
            .I(N__49592));
    LocalMux I__11105 (
            .O(N__49640),
            .I(N__49589));
    InMux I__11104 (
            .O(N__49639),
            .I(N__49586));
    InMux I__11103 (
            .O(N__49636),
            .I(N__49583));
    InMux I__11102 (
            .O(N__49635),
            .I(N__49572));
    InMux I__11101 (
            .O(N__49634),
            .I(N__49572));
    InMux I__11100 (
            .O(N__49631),
            .I(N__49572));
    InMux I__11099 (
            .O(N__49628),
            .I(N__49572));
    InMux I__11098 (
            .O(N__49625),
            .I(N__49572));
    InMux I__11097 (
            .O(N__49624),
            .I(N__49569));
    InMux I__11096 (
            .O(N__49623),
            .I(N__49564));
    InMux I__11095 (
            .O(N__49622),
            .I(N__49564));
    CascadeMux I__11094 (
            .O(N__49621),
            .I(N__49535));
    CascadeMux I__11093 (
            .O(N__49620),
            .I(N__49531));
    CascadeMux I__11092 (
            .O(N__49619),
            .I(N__49527));
    CascadeMux I__11091 (
            .O(N__49618),
            .I(N__49523));
    CascadeMux I__11090 (
            .O(N__49617),
            .I(N__49519));
    CascadeMux I__11089 (
            .O(N__49616),
            .I(N__49515));
    CascadeMux I__11088 (
            .O(N__49615),
            .I(N__49511));
    CascadeMux I__11087 (
            .O(N__49614),
            .I(N__49496));
    CascadeMux I__11086 (
            .O(N__49613),
            .I(N__49492));
    CascadeMux I__11085 (
            .O(N__49612),
            .I(N__49488));
    LocalMux I__11084 (
            .O(N__49609),
            .I(N__49484));
    Span4Mux_v I__11083 (
            .O(N__49606),
            .I(N__49477));
    Span4Mux_v I__11082 (
            .O(N__49597),
            .I(N__49477));
    LocalMux I__11081 (
            .O(N__49592),
            .I(N__49477));
    Span4Mux_v I__11080 (
            .O(N__49589),
            .I(N__49468));
    LocalMux I__11079 (
            .O(N__49586),
            .I(N__49468));
    LocalMux I__11078 (
            .O(N__49583),
            .I(N__49468));
    LocalMux I__11077 (
            .O(N__49572),
            .I(N__49468));
    LocalMux I__11076 (
            .O(N__49569),
            .I(N__49463));
    LocalMux I__11075 (
            .O(N__49564),
            .I(N__49463));
    InMux I__11074 (
            .O(N__49563),
            .I(N__49460));
    CascadeMux I__11073 (
            .O(N__49562),
            .I(N__49456));
    InMux I__11072 (
            .O(N__49561),
            .I(N__49441));
    InMux I__11071 (
            .O(N__49560),
            .I(N__49441));
    InMux I__11070 (
            .O(N__49559),
            .I(N__49441));
    InMux I__11069 (
            .O(N__49558),
            .I(N__49441));
    InMux I__11068 (
            .O(N__49557),
            .I(N__49441));
    InMux I__11067 (
            .O(N__49556),
            .I(N__49441));
    InMux I__11066 (
            .O(N__49555),
            .I(N__49441));
    InMux I__11065 (
            .O(N__49554),
            .I(N__49434));
    InMux I__11064 (
            .O(N__49553),
            .I(N__49434));
    InMux I__11063 (
            .O(N__49552),
            .I(N__49434));
    CascadeMux I__11062 (
            .O(N__49551),
            .I(N__49429));
    CascadeMux I__11061 (
            .O(N__49550),
            .I(N__49425));
    CascadeMux I__11060 (
            .O(N__49549),
            .I(N__49421));
    CascadeMux I__11059 (
            .O(N__49548),
            .I(N__49417));
    CascadeMux I__11058 (
            .O(N__49547),
            .I(N__49413));
    CascadeMux I__11057 (
            .O(N__49546),
            .I(N__49409));
    CascadeMux I__11056 (
            .O(N__49545),
            .I(N__49405));
    InMux I__11055 (
            .O(N__49544),
            .I(N__49399));
    InMux I__11054 (
            .O(N__49543),
            .I(N__49399));
    InMux I__11053 (
            .O(N__49542),
            .I(N__49390));
    InMux I__11052 (
            .O(N__49541),
            .I(N__49390));
    InMux I__11051 (
            .O(N__49540),
            .I(N__49390));
    InMux I__11050 (
            .O(N__49539),
            .I(N__49390));
    InMux I__11049 (
            .O(N__49538),
            .I(N__49375));
    InMux I__11048 (
            .O(N__49535),
            .I(N__49375));
    InMux I__11047 (
            .O(N__49534),
            .I(N__49375));
    InMux I__11046 (
            .O(N__49531),
            .I(N__49375));
    InMux I__11045 (
            .O(N__49530),
            .I(N__49375));
    InMux I__11044 (
            .O(N__49527),
            .I(N__49375));
    InMux I__11043 (
            .O(N__49526),
            .I(N__49375));
    InMux I__11042 (
            .O(N__49523),
            .I(N__49358));
    InMux I__11041 (
            .O(N__49522),
            .I(N__49358));
    InMux I__11040 (
            .O(N__49519),
            .I(N__49358));
    InMux I__11039 (
            .O(N__49518),
            .I(N__49358));
    InMux I__11038 (
            .O(N__49515),
            .I(N__49358));
    InMux I__11037 (
            .O(N__49514),
            .I(N__49358));
    InMux I__11036 (
            .O(N__49511),
            .I(N__49358));
    InMux I__11035 (
            .O(N__49510),
            .I(N__49358));
    CascadeMux I__11034 (
            .O(N__49509),
            .I(N__49355));
    CascadeMux I__11033 (
            .O(N__49508),
            .I(N__49351));
    CascadeMux I__11032 (
            .O(N__49507),
            .I(N__49347));
    CascadeMux I__11031 (
            .O(N__49506),
            .I(N__49343));
    CascadeMux I__11030 (
            .O(N__49505),
            .I(N__49339));
    CascadeMux I__11029 (
            .O(N__49504),
            .I(N__49335));
    CascadeMux I__11028 (
            .O(N__49503),
            .I(N__49331));
    CascadeMux I__11027 (
            .O(N__49502),
            .I(N__49327));
    CascadeMux I__11026 (
            .O(N__49501),
            .I(N__49323));
    CascadeMux I__11025 (
            .O(N__49500),
            .I(N__49319));
    CascadeMux I__11024 (
            .O(N__49499),
            .I(N__49315));
    InMux I__11023 (
            .O(N__49496),
            .I(N__49301));
    InMux I__11022 (
            .O(N__49495),
            .I(N__49301));
    InMux I__11021 (
            .O(N__49492),
            .I(N__49301));
    InMux I__11020 (
            .O(N__49491),
            .I(N__49301));
    InMux I__11019 (
            .O(N__49488),
            .I(N__49301));
    InMux I__11018 (
            .O(N__49487),
            .I(N__49301));
    Span12Mux_h I__11017 (
            .O(N__49484),
            .I(N__49298));
    Span4Mux_h I__11016 (
            .O(N__49477),
            .I(N__49295));
    Span4Mux_h I__11015 (
            .O(N__49468),
            .I(N__49292));
    Span4Mux_v I__11014 (
            .O(N__49463),
            .I(N__49287));
    LocalMux I__11013 (
            .O(N__49460),
            .I(N__49287));
    InMux I__11012 (
            .O(N__49459),
            .I(N__49282));
    InMux I__11011 (
            .O(N__49456),
            .I(N__49282));
    LocalMux I__11010 (
            .O(N__49441),
            .I(N__49277));
    LocalMux I__11009 (
            .O(N__49434),
            .I(N__49277));
    InMux I__11008 (
            .O(N__49433),
            .I(N__49260));
    InMux I__11007 (
            .O(N__49432),
            .I(N__49260));
    InMux I__11006 (
            .O(N__49429),
            .I(N__49260));
    InMux I__11005 (
            .O(N__49428),
            .I(N__49260));
    InMux I__11004 (
            .O(N__49425),
            .I(N__49260));
    InMux I__11003 (
            .O(N__49424),
            .I(N__49260));
    InMux I__11002 (
            .O(N__49421),
            .I(N__49260));
    InMux I__11001 (
            .O(N__49420),
            .I(N__49260));
    InMux I__11000 (
            .O(N__49417),
            .I(N__49243));
    InMux I__10999 (
            .O(N__49416),
            .I(N__49243));
    InMux I__10998 (
            .O(N__49413),
            .I(N__49243));
    InMux I__10997 (
            .O(N__49412),
            .I(N__49243));
    InMux I__10996 (
            .O(N__49409),
            .I(N__49243));
    InMux I__10995 (
            .O(N__49408),
            .I(N__49243));
    InMux I__10994 (
            .O(N__49405),
            .I(N__49243));
    InMux I__10993 (
            .O(N__49404),
            .I(N__49243));
    LocalMux I__10992 (
            .O(N__49399),
            .I(N__49234));
    LocalMux I__10991 (
            .O(N__49390),
            .I(N__49234));
    LocalMux I__10990 (
            .O(N__49375),
            .I(N__49234));
    LocalMux I__10989 (
            .O(N__49358),
            .I(N__49234));
    InMux I__10988 (
            .O(N__49355),
            .I(N__49217));
    InMux I__10987 (
            .O(N__49354),
            .I(N__49217));
    InMux I__10986 (
            .O(N__49351),
            .I(N__49217));
    InMux I__10985 (
            .O(N__49350),
            .I(N__49217));
    InMux I__10984 (
            .O(N__49347),
            .I(N__49217));
    InMux I__10983 (
            .O(N__49346),
            .I(N__49217));
    InMux I__10982 (
            .O(N__49343),
            .I(N__49217));
    InMux I__10981 (
            .O(N__49342),
            .I(N__49217));
    InMux I__10980 (
            .O(N__49339),
            .I(N__49200));
    InMux I__10979 (
            .O(N__49338),
            .I(N__49200));
    InMux I__10978 (
            .O(N__49335),
            .I(N__49200));
    InMux I__10977 (
            .O(N__49334),
            .I(N__49200));
    InMux I__10976 (
            .O(N__49331),
            .I(N__49200));
    InMux I__10975 (
            .O(N__49330),
            .I(N__49200));
    InMux I__10974 (
            .O(N__49327),
            .I(N__49200));
    InMux I__10973 (
            .O(N__49326),
            .I(N__49200));
    InMux I__10972 (
            .O(N__49323),
            .I(N__49187));
    InMux I__10971 (
            .O(N__49322),
            .I(N__49187));
    InMux I__10970 (
            .O(N__49319),
            .I(N__49187));
    InMux I__10969 (
            .O(N__49318),
            .I(N__49187));
    InMux I__10968 (
            .O(N__49315),
            .I(N__49187));
    InMux I__10967 (
            .O(N__49314),
            .I(N__49187));
    LocalMux I__10966 (
            .O(N__49301),
            .I(N__49184));
    Odrv12 I__10965 (
            .O(N__49298),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10964 (
            .O(N__49295),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10963 (
            .O(N__49292),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10962 (
            .O(N__49287),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10961 (
            .O(N__49282),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__10960 (
            .O(N__49277),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10959 (
            .O(N__49260),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10958 (
            .O(N__49243),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10957 (
            .O(N__49234),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10956 (
            .O(N__49217),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10955 (
            .O(N__49200),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10954 (
            .O(N__49187),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10953 (
            .O(N__49184),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__10952 (
            .O(N__49157),
            .I(N__49154));
    LocalMux I__10951 (
            .O(N__49154),
            .I(N__49151));
    Span4Mux_h I__10950 (
            .O(N__49151),
            .I(N__49148));
    Odrv4 I__10949 (
            .O(N__49148),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ));
    InMux I__10948 (
            .O(N__49145),
            .I(N__49138));
    InMux I__10947 (
            .O(N__49144),
            .I(N__49138));
    InMux I__10946 (
            .O(N__49143),
            .I(N__49135));
    LocalMux I__10945 (
            .O(N__49138),
            .I(N__49130));
    LocalMux I__10944 (
            .O(N__49135),
            .I(N__49130));
    Span4Mux_v I__10943 (
            .O(N__49130),
            .I(N__49125));
    CascadeMux I__10942 (
            .O(N__49129),
            .I(N__49122));
    CascadeMux I__10941 (
            .O(N__49128),
            .I(N__49119));
    Span4Mux_h I__10940 (
            .O(N__49125),
            .I(N__49115));
    InMux I__10939 (
            .O(N__49122),
            .I(N__49110));
    InMux I__10938 (
            .O(N__49119),
            .I(N__49110));
    InMux I__10937 (
            .O(N__49118),
            .I(N__49107));
    Span4Mux_h I__10936 (
            .O(N__49115),
            .I(N__49104));
    LocalMux I__10935 (
            .O(N__49110),
            .I(state_3));
    LocalMux I__10934 (
            .O(N__49107),
            .I(state_3));
    Odrv4 I__10933 (
            .O(N__49104),
            .I(state_3));
    IoInMux I__10932 (
            .O(N__49097),
            .I(N__49094));
    LocalMux I__10931 (
            .O(N__49094),
            .I(N__49091));
    Span4Mux_s2_v I__10930 (
            .O(N__49091),
            .I(N__49088));
    Span4Mux_v I__10929 (
            .O(N__49088),
            .I(N__49085));
    Span4Mux_v I__10928 (
            .O(N__49085),
            .I(N__49080));
    InMux I__10927 (
            .O(N__49084),
            .I(N__49075));
    InMux I__10926 (
            .O(N__49083),
            .I(N__49075));
    Span4Mux_v I__10925 (
            .O(N__49080),
            .I(N__49072));
    LocalMux I__10924 (
            .O(N__49075),
            .I(N__49069));
    Odrv4 I__10923 (
            .O(N__49072),
            .I(s1_phy_c));
    Odrv4 I__10922 (
            .O(N__49069),
            .I(s1_phy_c));
    InMux I__10921 (
            .O(N__49064),
            .I(N__49058));
    InMux I__10920 (
            .O(N__49063),
            .I(N__49055));
    InMux I__10919 (
            .O(N__49062),
            .I(N__49052));
    InMux I__10918 (
            .O(N__49061),
            .I(N__49049));
    LocalMux I__10917 (
            .O(N__49058),
            .I(N__49046));
    LocalMux I__10916 (
            .O(N__49055),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__10915 (
            .O(N__49052),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__10914 (
            .O(N__49049),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__10913 (
            .O(N__49046),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    CascadeMux I__10912 (
            .O(N__49037),
            .I(N__49033));
    InMux I__10911 (
            .O(N__49036),
            .I(N__49028));
    InMux I__10910 (
            .O(N__49033),
            .I(N__49023));
    InMux I__10909 (
            .O(N__49032),
            .I(N__49023));
    InMux I__10908 (
            .O(N__49031),
            .I(N__49020));
    LocalMux I__10907 (
            .O(N__49028),
            .I(N__49017));
    LocalMux I__10906 (
            .O(N__49023),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__10905 (
            .O(N__49020),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__10904 (
            .O(N__49017),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__10903 (
            .O(N__49010),
            .I(N__49007));
    LocalMux I__10902 (
            .O(N__49007),
            .I(N__49004));
    Span4Mux_s0_v I__10901 (
            .O(N__49004),
            .I(N__49001));
    Span4Mux_h I__10900 (
            .O(N__49001),
            .I(N__48998));
    Sp12to4 I__10899 (
            .O(N__48998),
            .I(N__48995));
    Span12Mux_v I__10898 (
            .O(N__48995),
            .I(N__48992));
    Odrv12 I__10897 (
            .O(N__48992),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    InMux I__10896 (
            .O(N__48989),
            .I(N__48986));
    LocalMux I__10895 (
            .O(N__48986),
            .I(N__48983));
    Span4Mux_s2_h I__10894 (
            .O(N__48983),
            .I(N__48979));
    InMux I__10893 (
            .O(N__48982),
            .I(N__48976));
    Span4Mux_h I__10892 (
            .O(N__48979),
            .I(N__48973));
    LocalMux I__10891 (
            .O(N__48976),
            .I(N__48968));
    Span4Mux_v I__10890 (
            .O(N__48973),
            .I(N__48968));
    Odrv4 I__10889 (
            .O(N__48968),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__10888 (
            .O(N__48965),
            .I(N__48961));
    InMux I__10887 (
            .O(N__48964),
            .I(N__48958));
    LocalMux I__10886 (
            .O(N__48961),
            .I(N__48955));
    LocalMux I__10885 (
            .O(N__48958),
            .I(N__48950));
    Span12Mux_s9_v I__10884 (
            .O(N__48955),
            .I(N__48950));
    Odrv12 I__10883 (
            .O(N__48950),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__10882 (
            .O(N__48947),
            .I(N__48944));
    LocalMux I__10881 (
            .O(N__48944),
            .I(N__48941));
    Span4Mux_s2_h I__10880 (
            .O(N__48941),
            .I(N__48937));
    InMux I__10879 (
            .O(N__48940),
            .I(N__48934));
    Span4Mux_h I__10878 (
            .O(N__48937),
            .I(N__48931));
    LocalMux I__10877 (
            .O(N__48934),
            .I(N__48926));
    Span4Mux_v I__10876 (
            .O(N__48931),
            .I(N__48926));
    Odrv4 I__10875 (
            .O(N__48926),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__10874 (
            .O(N__48923),
            .I(N__48920));
    LocalMux I__10873 (
            .O(N__48920),
            .I(N__48916));
    InMux I__10872 (
            .O(N__48919),
            .I(N__48913));
    Span4Mux_v I__10871 (
            .O(N__48916),
            .I(N__48910));
    LocalMux I__10870 (
            .O(N__48913),
            .I(N__48905));
    Span4Mux_h I__10869 (
            .O(N__48910),
            .I(N__48905));
    Span4Mux_h I__10868 (
            .O(N__48905),
            .I(N__48902));
    Odrv4 I__10867 (
            .O(N__48902),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    CascadeMux I__10866 (
            .O(N__48899),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_cascade_ ));
    InMux I__10865 (
            .O(N__48896),
            .I(N__48893));
    LocalMux I__10864 (
            .O(N__48893),
            .I(N__48890));
    Span4Mux_s3_v I__10863 (
            .O(N__48890),
            .I(N__48887));
    Odrv4 I__10862 (
            .O(N__48887),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__10861 (
            .O(N__48884),
            .I(N__48881));
    LocalMux I__10860 (
            .O(N__48881),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__10859 (
            .O(N__48878),
            .I(N__48872));
    InMux I__10858 (
            .O(N__48877),
            .I(N__48872));
    LocalMux I__10857 (
            .O(N__48872),
            .I(N__48867));
    InMux I__10856 (
            .O(N__48871),
            .I(N__48862));
    InMux I__10855 (
            .O(N__48870),
            .I(N__48862));
    Span4Mux_h I__10854 (
            .O(N__48867),
            .I(N__48859));
    LocalMux I__10853 (
            .O(N__48862),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__10852 (
            .O(N__48859),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    CascadeMux I__10851 (
            .O(N__48854),
            .I(N__48850));
    InMux I__10850 (
            .O(N__48853),
            .I(N__48842));
    InMux I__10849 (
            .O(N__48850),
            .I(N__48842));
    InMux I__10848 (
            .O(N__48849),
            .I(N__48842));
    LocalMux I__10847 (
            .O(N__48842),
            .I(N__48839));
    Span4Mux_h I__10846 (
            .O(N__48839),
            .I(N__48836));
    Odrv4 I__10845 (
            .O(N__48836),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    ClkMux I__10844 (
            .O(N__48833),
            .I(N__48830));
    GlobalMux I__10843 (
            .O(N__48830),
            .I(N__48827));
    gio2CtrlBuf I__10842 (
            .O(N__48827),
            .I(delay_tr_input_c_g));
    CEMux I__10841 (
            .O(N__48824),
            .I(N__48821));
    LocalMux I__10840 (
            .O(N__48821),
            .I(N__48818));
    Span4Mux_v I__10839 (
            .O(N__48818),
            .I(N__48812));
    CEMux I__10838 (
            .O(N__48817),
            .I(N__48809));
    CEMux I__10837 (
            .O(N__48816),
            .I(N__48806));
    CEMux I__10836 (
            .O(N__48815),
            .I(N__48803));
    Odrv4 I__10835 (
            .O(N__48812),
            .I(\current_shift_inst.timer_s1.N_164_i ));
    LocalMux I__10834 (
            .O(N__48809),
            .I(\current_shift_inst.timer_s1.N_164_i ));
    LocalMux I__10833 (
            .O(N__48806),
            .I(\current_shift_inst.timer_s1.N_164_i ));
    LocalMux I__10832 (
            .O(N__48803),
            .I(\current_shift_inst.timer_s1.N_164_i ));
    InMux I__10831 (
            .O(N__48794),
            .I(N__48784));
    InMux I__10830 (
            .O(N__48793),
            .I(N__48784));
    InMux I__10829 (
            .O(N__48792),
            .I(N__48784));
    InMux I__10828 (
            .O(N__48791),
            .I(N__48781));
    LocalMux I__10827 (
            .O(N__48784),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__10826 (
            .O(N__48781),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__10825 (
            .O(N__48776),
            .I(N__48756));
    InMux I__10824 (
            .O(N__48775),
            .I(N__48756));
    InMux I__10823 (
            .O(N__48774),
            .I(N__48756));
    InMux I__10822 (
            .O(N__48773),
            .I(N__48756));
    InMux I__10821 (
            .O(N__48772),
            .I(N__48735));
    InMux I__10820 (
            .O(N__48771),
            .I(N__48735));
    InMux I__10819 (
            .O(N__48770),
            .I(N__48735));
    InMux I__10818 (
            .O(N__48769),
            .I(N__48735));
    InMux I__10817 (
            .O(N__48768),
            .I(N__48726));
    InMux I__10816 (
            .O(N__48767),
            .I(N__48726));
    InMux I__10815 (
            .O(N__48766),
            .I(N__48726));
    InMux I__10814 (
            .O(N__48765),
            .I(N__48726));
    LocalMux I__10813 (
            .O(N__48756),
            .I(N__48717));
    InMux I__10812 (
            .O(N__48755),
            .I(N__48708));
    InMux I__10811 (
            .O(N__48754),
            .I(N__48708));
    InMux I__10810 (
            .O(N__48753),
            .I(N__48708));
    InMux I__10809 (
            .O(N__48752),
            .I(N__48708));
    InMux I__10808 (
            .O(N__48751),
            .I(N__48699));
    InMux I__10807 (
            .O(N__48750),
            .I(N__48699));
    InMux I__10806 (
            .O(N__48749),
            .I(N__48699));
    InMux I__10805 (
            .O(N__48748),
            .I(N__48699));
    InMux I__10804 (
            .O(N__48747),
            .I(N__48690));
    InMux I__10803 (
            .O(N__48746),
            .I(N__48690));
    InMux I__10802 (
            .O(N__48745),
            .I(N__48690));
    InMux I__10801 (
            .O(N__48744),
            .I(N__48690));
    LocalMux I__10800 (
            .O(N__48735),
            .I(N__48685));
    LocalMux I__10799 (
            .O(N__48726),
            .I(N__48685));
    InMux I__10798 (
            .O(N__48725),
            .I(N__48680));
    InMux I__10797 (
            .O(N__48724),
            .I(N__48680));
    InMux I__10796 (
            .O(N__48723),
            .I(N__48671));
    InMux I__10795 (
            .O(N__48722),
            .I(N__48671));
    InMux I__10794 (
            .O(N__48721),
            .I(N__48671));
    InMux I__10793 (
            .O(N__48720),
            .I(N__48671));
    Span4Mux_h I__10792 (
            .O(N__48717),
            .I(N__48668));
    LocalMux I__10791 (
            .O(N__48708),
            .I(N__48659));
    LocalMux I__10790 (
            .O(N__48699),
            .I(N__48659));
    LocalMux I__10789 (
            .O(N__48690),
            .I(N__48659));
    Span4Mux_h I__10788 (
            .O(N__48685),
            .I(N__48659));
    LocalMux I__10787 (
            .O(N__48680),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__10786 (
            .O(N__48671),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__10785 (
            .O(N__48668),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__10784 (
            .O(N__48659),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__10783 (
            .O(N__48650),
            .I(N__48647));
    LocalMux I__10782 (
            .O(N__48647),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ));
    InMux I__10781 (
            .O(N__48644),
            .I(N__48641));
    LocalMux I__10780 (
            .O(N__48641),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    CascadeMux I__10779 (
            .O(N__48638),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ));
    InMux I__10778 (
            .O(N__48635),
            .I(N__48632));
    LocalMux I__10777 (
            .O(N__48632),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    InMux I__10776 (
            .O(N__48629),
            .I(N__48626));
    LocalMux I__10775 (
            .O(N__48626),
            .I(N__48623));
    Odrv4 I__10774 (
            .O(N__48623),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    CascadeMux I__10773 (
            .O(N__48620),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ));
    InMux I__10772 (
            .O(N__48617),
            .I(N__48614));
    LocalMux I__10771 (
            .O(N__48614),
            .I(N__48611));
    Odrv12 I__10770 (
            .O(N__48611),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__10769 (
            .O(N__48608),
            .I(N__48605));
    LocalMux I__10768 (
            .O(N__48605),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ));
    InMux I__10767 (
            .O(N__48602),
            .I(N__48599));
    LocalMux I__10766 (
            .O(N__48599),
            .I(N__48596));
    Odrv4 I__10765 (
            .O(N__48596),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__10764 (
            .O(N__48593),
            .I(N__48590));
    LocalMux I__10763 (
            .O(N__48590),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    CascadeMux I__10762 (
            .O(N__48587),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ));
    CascadeMux I__10761 (
            .O(N__48584),
            .I(\current_shift_inst.PI_CTRL.N_47_cascade_ ));
    InMux I__10760 (
            .O(N__48581),
            .I(N__48578));
    LocalMux I__10759 (
            .O(N__48578),
            .I(\current_shift_inst.PI_CTRL.N_46_21 ));
    CascadeMux I__10758 (
            .O(N__48575),
            .I(N__48572));
    InMux I__10757 (
            .O(N__48572),
            .I(N__48569));
    LocalMux I__10756 (
            .O(N__48569),
            .I(N__48566));
    Span4Mux_v I__10755 (
            .O(N__48566),
            .I(N__48563));
    Span4Mux_h I__10754 (
            .O(N__48563),
            .I(N__48560));
    Odrv4 I__10753 (
            .O(N__48560),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__10752 (
            .O(N__48557),
            .I(N__48554));
    LocalMux I__10751 (
            .O(N__48554),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__10750 (
            .O(N__48551),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    InMux I__10749 (
            .O(N__48548),
            .I(N__48545));
    LocalMux I__10748 (
            .O(N__48545),
            .I(N__48542));
    Span12Mux_s6_v I__10747 (
            .O(N__48542),
            .I(N__48539));
    Odrv12 I__10746 (
            .O(N__48539),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__10745 (
            .O(N__48536),
            .I(N__48533));
    LocalMux I__10744 (
            .O(N__48533),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__10743 (
            .O(N__48530),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    InMux I__10742 (
            .O(N__48527),
            .I(N__48524));
    LocalMux I__10741 (
            .O(N__48524),
            .I(N__48521));
    Span4Mux_h I__10740 (
            .O(N__48521),
            .I(N__48518));
    Span4Mux_h I__10739 (
            .O(N__48518),
            .I(N__48515));
    Odrv4 I__10738 (
            .O(N__48515),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__10737 (
            .O(N__48512),
            .I(N__48509));
    LocalMux I__10736 (
            .O(N__48509),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__10735 (
            .O(N__48506),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__10734 (
            .O(N__48503),
            .I(N__48500));
    InMux I__10733 (
            .O(N__48500),
            .I(N__48497));
    LocalMux I__10732 (
            .O(N__48497),
            .I(N__48494));
    Span4Mux_h I__10731 (
            .O(N__48494),
            .I(N__48491));
    Span4Mux_h I__10730 (
            .O(N__48491),
            .I(N__48488));
    Odrv4 I__10729 (
            .O(N__48488),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__10728 (
            .O(N__48485),
            .I(N__48482));
    LocalMux I__10727 (
            .O(N__48482),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__10726 (
            .O(N__48479),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    InMux I__10725 (
            .O(N__48476),
            .I(N__48473));
    LocalMux I__10724 (
            .O(N__48473),
            .I(N__48470));
    Span4Mux_h I__10723 (
            .O(N__48470),
            .I(N__48467));
    Span4Mux_h I__10722 (
            .O(N__48467),
            .I(N__48464));
    Odrv4 I__10721 (
            .O(N__48464),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__10720 (
            .O(N__48461),
            .I(N__48458));
    LocalMux I__10719 (
            .O(N__48458),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__10718 (
            .O(N__48455),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__10717 (
            .O(N__48452),
            .I(N__48449));
    LocalMux I__10716 (
            .O(N__48449),
            .I(N__48446));
    Span4Mux_v I__10715 (
            .O(N__48446),
            .I(N__48443));
    Span4Mux_h I__10714 (
            .O(N__48443),
            .I(N__48440));
    Odrv4 I__10713 (
            .O(N__48440),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30 ));
    CascadeMux I__10712 (
            .O(N__48437),
            .I(N__48434));
    InMux I__10711 (
            .O(N__48434),
            .I(N__48431));
    LocalMux I__10710 (
            .O(N__48431),
            .I(N__48428));
    Span4Mux_h I__10709 (
            .O(N__48428),
            .I(N__48425));
    Span4Mux_h I__10708 (
            .O(N__48425),
            .I(N__48422));
    Odrv4 I__10707 (
            .O(N__48422),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    InMux I__10706 (
            .O(N__48419),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    CascadeMux I__10705 (
            .O(N__48416),
            .I(N__48413));
    InMux I__10704 (
            .O(N__48413),
            .I(N__48410));
    LocalMux I__10703 (
            .O(N__48410),
            .I(N__48407));
    Span4Mux_v I__10702 (
            .O(N__48407),
            .I(N__48404));
    Span4Mux_h I__10701 (
            .O(N__48404),
            .I(N__48401));
    Odrv4 I__10700 (
            .O(N__48401),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__10699 (
            .O(N__48398),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__10698 (
            .O(N__48395),
            .I(N__48392));
    InMux I__10697 (
            .O(N__48392),
            .I(N__48389));
    LocalMux I__10696 (
            .O(N__48389),
            .I(N__48386));
    Span4Mux_v I__10695 (
            .O(N__48386),
            .I(N__48383));
    Span4Mux_h I__10694 (
            .O(N__48383),
            .I(N__48380));
    Odrv4 I__10693 (
            .O(N__48380),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__10692 (
            .O(N__48377),
            .I(N__48374));
    LocalMux I__10691 (
            .O(N__48374),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__10690 (
            .O(N__48371),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    CascadeMux I__10689 (
            .O(N__48368),
            .I(N__48365));
    InMux I__10688 (
            .O(N__48365),
            .I(N__48362));
    LocalMux I__10687 (
            .O(N__48362),
            .I(N__48359));
    Span4Mux_h I__10686 (
            .O(N__48359),
            .I(N__48356));
    Span4Mux_h I__10685 (
            .O(N__48356),
            .I(N__48353));
    Odrv4 I__10684 (
            .O(N__48353),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__10683 (
            .O(N__48350),
            .I(N__48347));
    LocalMux I__10682 (
            .O(N__48347),
            .I(N__48344));
    Span4Mux_h I__10681 (
            .O(N__48344),
            .I(N__48341));
    Odrv4 I__10680 (
            .O(N__48341),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__10679 (
            .O(N__48338),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__10678 (
            .O(N__48335),
            .I(N__48332));
    InMux I__10677 (
            .O(N__48332),
            .I(N__48329));
    LocalMux I__10676 (
            .O(N__48329),
            .I(N__48326));
    Span4Mux_h I__10675 (
            .O(N__48326),
            .I(N__48323));
    Span4Mux_h I__10674 (
            .O(N__48323),
            .I(N__48320));
    Odrv4 I__10673 (
            .O(N__48320),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__10672 (
            .O(N__48317),
            .I(N__48314));
    LocalMux I__10671 (
            .O(N__48314),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__10670 (
            .O(N__48311),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__10669 (
            .O(N__48308),
            .I(N__48305));
    InMux I__10668 (
            .O(N__48305),
            .I(N__48302));
    LocalMux I__10667 (
            .O(N__48302),
            .I(N__48299));
    Span4Mux_h I__10666 (
            .O(N__48299),
            .I(N__48296));
    Span4Mux_h I__10665 (
            .O(N__48296),
            .I(N__48293));
    Odrv4 I__10664 (
            .O(N__48293),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__10663 (
            .O(N__48290),
            .I(N__48287));
    LocalMux I__10662 (
            .O(N__48287),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__10661 (
            .O(N__48284),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__10660 (
            .O(N__48281),
            .I(N__48278));
    InMux I__10659 (
            .O(N__48278),
            .I(N__48275));
    LocalMux I__10658 (
            .O(N__48275),
            .I(N__48272));
    Span4Mux_h I__10657 (
            .O(N__48272),
            .I(N__48269));
    Span4Mux_h I__10656 (
            .O(N__48269),
            .I(N__48266));
    Odrv4 I__10655 (
            .O(N__48266),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__10654 (
            .O(N__48263),
            .I(N__48260));
    LocalMux I__10653 (
            .O(N__48260),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__10652 (
            .O(N__48257),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    InMux I__10651 (
            .O(N__48254),
            .I(N__48251));
    LocalMux I__10650 (
            .O(N__48251),
            .I(N__48248));
    Span4Mux_h I__10649 (
            .O(N__48248),
            .I(N__48245));
    Span4Mux_h I__10648 (
            .O(N__48245),
            .I(N__48242));
    Odrv4 I__10647 (
            .O(N__48242),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__10646 (
            .O(N__48239),
            .I(N__48236));
    LocalMux I__10645 (
            .O(N__48236),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__10644 (
            .O(N__48233),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    InMux I__10643 (
            .O(N__48230),
            .I(N__48227));
    LocalMux I__10642 (
            .O(N__48227),
            .I(N__48224));
    Span4Mux_h I__10641 (
            .O(N__48224),
            .I(N__48221));
    Span4Mux_h I__10640 (
            .O(N__48221),
            .I(N__48218));
    Odrv4 I__10639 (
            .O(N__48218),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__10638 (
            .O(N__48215),
            .I(N__48212));
    LocalMux I__10637 (
            .O(N__48212),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__10636 (
            .O(N__48209),
            .I(bfn_17_26_0_));
    CascadeMux I__10635 (
            .O(N__48206),
            .I(N__48203));
    InMux I__10634 (
            .O(N__48203),
            .I(N__48200));
    LocalMux I__10633 (
            .O(N__48200),
            .I(N__48197));
    Span4Mux_h I__10632 (
            .O(N__48197),
            .I(N__48194));
    Span4Mux_h I__10631 (
            .O(N__48194),
            .I(N__48191));
    Odrv4 I__10630 (
            .O(N__48191),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__10629 (
            .O(N__48188),
            .I(N__48185));
    LocalMux I__10628 (
            .O(N__48185),
            .I(N__48182));
    Span4Mux_v I__10627 (
            .O(N__48182),
            .I(N__48179));
    Odrv4 I__10626 (
            .O(N__48179),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__10625 (
            .O(N__48176),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__10624 (
            .O(N__48173),
            .I(N__48170));
    InMux I__10623 (
            .O(N__48170),
            .I(N__48167));
    LocalMux I__10622 (
            .O(N__48167),
            .I(N__48164));
    Span4Mux_h I__10621 (
            .O(N__48164),
            .I(N__48161));
    Span4Mux_h I__10620 (
            .O(N__48161),
            .I(N__48158));
    Odrv4 I__10619 (
            .O(N__48158),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__10618 (
            .O(N__48155),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    CascadeMux I__10617 (
            .O(N__48152),
            .I(N__48149));
    InMux I__10616 (
            .O(N__48149),
            .I(N__48146));
    LocalMux I__10615 (
            .O(N__48146),
            .I(N__48143));
    Span4Mux_h I__10614 (
            .O(N__48143),
            .I(N__48140));
    Span4Mux_h I__10613 (
            .O(N__48140),
            .I(N__48137));
    Odrv4 I__10612 (
            .O(N__48137),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__10611 (
            .O(N__48134),
            .I(N__48131));
    LocalMux I__10610 (
            .O(N__48131),
            .I(N__48128));
    Span4Mux_v I__10609 (
            .O(N__48128),
            .I(N__48125));
    Odrv4 I__10608 (
            .O(N__48125),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__10607 (
            .O(N__48122),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__10606 (
            .O(N__48119),
            .I(N__48116));
    InMux I__10605 (
            .O(N__48116),
            .I(N__48113));
    LocalMux I__10604 (
            .O(N__48113),
            .I(N__48110));
    Sp12to4 I__10603 (
            .O(N__48110),
            .I(N__48107));
    Odrv12 I__10602 (
            .O(N__48107),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__10601 (
            .O(N__48104),
            .I(N__48101));
    LocalMux I__10600 (
            .O(N__48101),
            .I(N__48098));
    Span4Mux_s3_v I__10599 (
            .O(N__48098),
            .I(N__48095));
    Odrv4 I__10598 (
            .O(N__48095),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__10597 (
            .O(N__48092),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    CascadeMux I__10596 (
            .O(N__48089),
            .I(N__48086));
    InMux I__10595 (
            .O(N__48086),
            .I(N__48083));
    LocalMux I__10594 (
            .O(N__48083),
            .I(N__48080));
    Odrv12 I__10593 (
            .O(N__48080),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__10592 (
            .O(N__48077),
            .I(N__48074));
    LocalMux I__10591 (
            .O(N__48074),
            .I(N__48071));
    Span4Mux_v I__10590 (
            .O(N__48071),
            .I(N__48068));
    Odrv4 I__10589 (
            .O(N__48068),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__10588 (
            .O(N__48065),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__10587 (
            .O(N__48062),
            .I(N__48059));
    InMux I__10586 (
            .O(N__48059),
            .I(N__48056));
    LocalMux I__10585 (
            .O(N__48056),
            .I(N__48053));
    Sp12to4 I__10584 (
            .O(N__48053),
            .I(N__48050));
    Odrv12 I__10583 (
            .O(N__48050),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__10582 (
            .O(N__48047),
            .I(N__48044));
    LocalMux I__10581 (
            .O(N__48044),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__10580 (
            .O(N__48041),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__10579 (
            .O(N__48038),
            .I(N__48035));
    InMux I__10578 (
            .O(N__48035),
            .I(N__48032));
    LocalMux I__10577 (
            .O(N__48032),
            .I(N__48029));
    Span4Mux_v I__10576 (
            .O(N__48029),
            .I(N__48026));
    Span4Mux_h I__10575 (
            .O(N__48026),
            .I(N__48023));
    Odrv4 I__10574 (
            .O(N__48023),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__10573 (
            .O(N__48020),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    CascadeMux I__10572 (
            .O(N__48017),
            .I(N__48014));
    InMux I__10571 (
            .O(N__48014),
            .I(N__48011));
    LocalMux I__10570 (
            .O(N__48011),
            .I(N__48008));
    Span4Mux_h I__10569 (
            .O(N__48008),
            .I(N__48005));
    Span4Mux_h I__10568 (
            .O(N__48005),
            .I(N__48002));
    Odrv4 I__10567 (
            .O(N__48002),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__10566 (
            .O(N__47999),
            .I(bfn_17_25_0_));
    CascadeMux I__10565 (
            .O(N__47996),
            .I(N__47993));
    InMux I__10564 (
            .O(N__47993),
            .I(N__47990));
    LocalMux I__10563 (
            .O(N__47990),
            .I(N__47987));
    Span4Mux_h I__10562 (
            .O(N__47987),
            .I(N__47984));
    Span4Mux_h I__10561 (
            .O(N__47984),
            .I(N__47981));
    Odrv4 I__10560 (
            .O(N__47981),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__10559 (
            .O(N__47978),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    CascadeMux I__10558 (
            .O(N__47975),
            .I(N__47972));
    InMux I__10557 (
            .O(N__47972),
            .I(N__47969));
    LocalMux I__10556 (
            .O(N__47969),
            .I(N__47966));
    Span4Mux_h I__10555 (
            .O(N__47966),
            .I(N__47963));
    Span4Mux_h I__10554 (
            .O(N__47963),
            .I(N__47960));
    Odrv4 I__10553 (
            .O(N__47960),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__10552 (
            .O(N__47957),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__10551 (
            .O(N__47954),
            .I(N__47951));
    InMux I__10550 (
            .O(N__47951),
            .I(N__47948));
    LocalMux I__10549 (
            .O(N__47948),
            .I(N__47945));
    Span4Mux_h I__10548 (
            .O(N__47945),
            .I(N__47942));
    Span4Mux_h I__10547 (
            .O(N__47942),
            .I(N__47939));
    Odrv4 I__10546 (
            .O(N__47939),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    InMux I__10545 (
            .O(N__47936),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__10544 (
            .O(N__47933),
            .I(N__47930));
    InMux I__10543 (
            .O(N__47930),
            .I(N__47927));
    LocalMux I__10542 (
            .O(N__47927),
            .I(N__47924));
    Span12Mux_v I__10541 (
            .O(N__47924),
            .I(N__47921));
    Odrv12 I__10540 (
            .O(N__47921),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__10539 (
            .O(N__47918),
            .I(N__47915));
    LocalMux I__10538 (
            .O(N__47915),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__10537 (
            .O(N__47912),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__10536 (
            .O(N__47909),
            .I(N__47906));
    InMux I__10535 (
            .O(N__47906),
            .I(N__47903));
    LocalMux I__10534 (
            .O(N__47903),
            .I(N__47900));
    Odrv12 I__10533 (
            .O(N__47900),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__10532 (
            .O(N__47897),
            .I(N__47894));
    LocalMux I__10531 (
            .O(N__47894),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__10530 (
            .O(N__47891),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__10529 (
            .O(N__47888),
            .I(N__47885));
    InMux I__10528 (
            .O(N__47885),
            .I(N__47882));
    LocalMux I__10527 (
            .O(N__47882),
            .I(N__47879));
    Span12Mux_h I__10526 (
            .O(N__47879),
            .I(N__47876));
    Odrv12 I__10525 (
            .O(N__47876),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__10524 (
            .O(N__47873),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__10523 (
            .O(N__47870),
            .I(N__47867));
    InMux I__10522 (
            .O(N__47867),
            .I(N__47864));
    LocalMux I__10521 (
            .O(N__47864),
            .I(N__47861));
    Odrv12 I__10520 (
            .O(N__47861),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__10519 (
            .O(N__47858),
            .I(N__47855));
    LocalMux I__10518 (
            .O(N__47855),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__10517 (
            .O(N__47852),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    InMux I__10516 (
            .O(N__47849),
            .I(N__47846));
    LocalMux I__10515 (
            .O(N__47846),
            .I(N__47843));
    Span4Mux_h I__10514 (
            .O(N__47843),
            .I(N__47840));
    Span4Mux_h I__10513 (
            .O(N__47840),
            .I(N__47837));
    Odrv4 I__10512 (
            .O(N__47837),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__10511 (
            .O(N__47834),
            .I(bfn_17_24_0_));
    InMux I__10510 (
            .O(N__47831),
            .I(N__47828));
    LocalMux I__10509 (
            .O(N__47828),
            .I(N__47825));
    Span4Mux_h I__10508 (
            .O(N__47825),
            .I(N__47822));
    Odrv4 I__10507 (
            .O(N__47822),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__10506 (
            .O(N__47819),
            .I(bfn_17_22_0_));
    InMux I__10505 (
            .O(N__47816),
            .I(N__47813));
    LocalMux I__10504 (
            .O(N__47813),
            .I(\current_shift_inst.control_input_axb_25 ));
    InMux I__10503 (
            .O(N__47810),
            .I(N__47807));
    LocalMux I__10502 (
            .O(N__47807),
            .I(N__47804));
    Span4Mux_h I__10501 (
            .O(N__47804),
            .I(N__47801));
    Odrv4 I__10500 (
            .O(N__47801),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__10499 (
            .O(N__47798),
            .I(\current_shift_inst.control_input_cry_24 ));
    InMux I__10498 (
            .O(N__47795),
            .I(N__47792));
    LocalMux I__10497 (
            .O(N__47792),
            .I(N__47789));
    Span4Mux_v I__10496 (
            .O(N__47789),
            .I(N__47786));
    Odrv4 I__10495 (
            .O(N__47786),
            .I(\current_shift_inst.control_input_axb_26 ));
    InMux I__10494 (
            .O(N__47783),
            .I(N__47780));
    LocalMux I__10493 (
            .O(N__47780),
            .I(N__47777));
    Span4Mux_v I__10492 (
            .O(N__47777),
            .I(N__47774));
    Odrv4 I__10491 (
            .O(N__47774),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ));
    InMux I__10490 (
            .O(N__47771),
            .I(\current_shift_inst.control_input_cry_25 ));
    InMux I__10489 (
            .O(N__47768),
            .I(N__47765));
    LocalMux I__10488 (
            .O(N__47765),
            .I(\current_shift_inst.control_input_axb_27 ));
    InMux I__10487 (
            .O(N__47762),
            .I(N__47759));
    LocalMux I__10486 (
            .O(N__47759),
            .I(N__47756));
    Span4Mux_v I__10485 (
            .O(N__47756),
            .I(N__47753));
    Odrv4 I__10484 (
            .O(N__47753),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ));
    InMux I__10483 (
            .O(N__47750),
            .I(\current_shift_inst.control_input_cry_26 ));
    InMux I__10482 (
            .O(N__47747),
            .I(N__47744));
    LocalMux I__10481 (
            .O(N__47744),
            .I(N__47741));
    Odrv12 I__10480 (
            .O(N__47741),
            .I(\current_shift_inst.control_input_axb_28 ));
    InMux I__10479 (
            .O(N__47738),
            .I(N__47735));
    LocalMux I__10478 (
            .O(N__47735),
            .I(N__47732));
    Span4Mux_h I__10477 (
            .O(N__47732),
            .I(N__47729));
    Odrv4 I__10476 (
            .O(N__47729),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ));
    InMux I__10475 (
            .O(N__47726),
            .I(\current_shift_inst.control_input_cry_27 ));
    InMux I__10474 (
            .O(N__47723),
            .I(N__47720));
    LocalMux I__10473 (
            .O(N__47720),
            .I(N__47717));
    Span4Mux_h I__10472 (
            .O(N__47717),
            .I(N__47714));
    Odrv4 I__10471 (
            .O(N__47714),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ));
    InMux I__10470 (
            .O(N__47711),
            .I(\current_shift_inst.control_input_cry_28 ));
    InMux I__10469 (
            .O(N__47708),
            .I(\current_shift_inst.control_input_cry_29 ));
    InMux I__10468 (
            .O(N__47705),
            .I(N__47702));
    LocalMux I__10467 (
            .O(N__47702),
            .I(N__47699));
    Span4Mux_h I__10466 (
            .O(N__47699),
            .I(N__47695));
    InMux I__10465 (
            .O(N__47698),
            .I(N__47692));
    Odrv4 I__10464 (
            .O(N__47695),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__10463 (
            .O(N__47692),
            .I(\current_shift_inst.control_input_31 ));
    CascadeMux I__10462 (
            .O(N__47687),
            .I(N__47682));
    InMux I__10461 (
            .O(N__47686),
            .I(N__47675));
    InMux I__10460 (
            .O(N__47685),
            .I(N__47675));
    InMux I__10459 (
            .O(N__47682),
            .I(N__47672));
    InMux I__10458 (
            .O(N__47681),
            .I(N__47666));
    InMux I__10457 (
            .O(N__47680),
            .I(N__47666));
    LocalMux I__10456 (
            .O(N__47675),
            .I(N__47656));
    LocalMux I__10455 (
            .O(N__47672),
            .I(N__47653));
    InMux I__10454 (
            .O(N__47671),
            .I(N__47644));
    LocalMux I__10453 (
            .O(N__47666),
            .I(N__47641));
    InMux I__10452 (
            .O(N__47665),
            .I(N__47636));
    InMux I__10451 (
            .O(N__47664),
            .I(N__47636));
    InMux I__10450 (
            .O(N__47663),
            .I(N__47625));
    InMux I__10449 (
            .O(N__47662),
            .I(N__47625));
    InMux I__10448 (
            .O(N__47661),
            .I(N__47625));
    InMux I__10447 (
            .O(N__47660),
            .I(N__47625));
    InMux I__10446 (
            .O(N__47659),
            .I(N__47625));
    Span4Mux_h I__10445 (
            .O(N__47656),
            .I(N__47609));
    Span4Mux_h I__10444 (
            .O(N__47653),
            .I(N__47606));
    InMux I__10443 (
            .O(N__47652),
            .I(N__47593));
    InMux I__10442 (
            .O(N__47651),
            .I(N__47593));
    InMux I__10441 (
            .O(N__47650),
            .I(N__47593));
    InMux I__10440 (
            .O(N__47649),
            .I(N__47593));
    InMux I__10439 (
            .O(N__47648),
            .I(N__47593));
    InMux I__10438 (
            .O(N__47647),
            .I(N__47593));
    LocalMux I__10437 (
            .O(N__47644),
            .I(N__47584));
    Span4Mux_h I__10436 (
            .O(N__47641),
            .I(N__47584));
    LocalMux I__10435 (
            .O(N__47636),
            .I(N__47584));
    LocalMux I__10434 (
            .O(N__47625),
            .I(N__47584));
    InMux I__10433 (
            .O(N__47624),
            .I(N__47567));
    InMux I__10432 (
            .O(N__47623),
            .I(N__47567));
    InMux I__10431 (
            .O(N__47622),
            .I(N__47567));
    InMux I__10430 (
            .O(N__47621),
            .I(N__47567));
    InMux I__10429 (
            .O(N__47620),
            .I(N__47567));
    InMux I__10428 (
            .O(N__47619),
            .I(N__47567));
    InMux I__10427 (
            .O(N__47618),
            .I(N__47567));
    InMux I__10426 (
            .O(N__47617),
            .I(N__47567));
    InMux I__10425 (
            .O(N__47616),
            .I(N__47556));
    InMux I__10424 (
            .O(N__47615),
            .I(N__47556));
    InMux I__10423 (
            .O(N__47614),
            .I(N__47556));
    InMux I__10422 (
            .O(N__47613),
            .I(N__47556));
    InMux I__10421 (
            .O(N__47612),
            .I(N__47556));
    Odrv4 I__10420 (
            .O(N__47609),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__10419 (
            .O(N__47606),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__10418 (
            .O(N__47593),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__10417 (
            .O(N__47584),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__10416 (
            .O(N__47567),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__10415 (
            .O(N__47556),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__10414 (
            .O(N__47543),
            .I(N__47540));
    LocalMux I__10413 (
            .O(N__47540),
            .I(\current_shift_inst.control_input_axb_29 ));
    CascadeMux I__10412 (
            .O(N__47537),
            .I(N__47534));
    InMux I__10411 (
            .O(N__47534),
            .I(N__47531));
    LocalMux I__10410 (
            .O(N__47531),
            .I(N__47528));
    Span4Mux_h I__10409 (
            .O(N__47528),
            .I(N__47525));
    Span4Mux_h I__10408 (
            .O(N__47525),
            .I(N__47522));
    Odrv4 I__10407 (
            .O(N__47522),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    InMux I__10406 (
            .O(N__47519),
            .I(N__47516));
    LocalMux I__10405 (
            .O(N__47516),
            .I(\current_shift_inst.control_input_axb_17 ));
    InMux I__10404 (
            .O(N__47513),
            .I(N__47510));
    LocalMux I__10403 (
            .O(N__47510),
            .I(N__47507));
    Span4Mux_h I__10402 (
            .O(N__47507),
            .I(N__47504));
    Odrv4 I__10401 (
            .O(N__47504),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__10400 (
            .O(N__47501),
            .I(\current_shift_inst.control_input_cry_16 ));
    InMux I__10399 (
            .O(N__47498),
            .I(N__47495));
    LocalMux I__10398 (
            .O(N__47495),
            .I(N__47492));
    Span4Mux_v I__10397 (
            .O(N__47492),
            .I(N__47489));
    Odrv4 I__10396 (
            .O(N__47489),
            .I(\current_shift_inst.control_input_axb_18 ));
    InMux I__10395 (
            .O(N__47486),
            .I(N__47483));
    LocalMux I__10394 (
            .O(N__47483),
            .I(N__47480));
    Span4Mux_v I__10393 (
            .O(N__47480),
            .I(N__47477));
    Odrv4 I__10392 (
            .O(N__47477),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    InMux I__10391 (
            .O(N__47474),
            .I(\current_shift_inst.control_input_cry_17 ));
    InMux I__10390 (
            .O(N__47471),
            .I(N__47468));
    LocalMux I__10389 (
            .O(N__47468),
            .I(N__47465));
    Span4Mux_v I__10388 (
            .O(N__47465),
            .I(N__47462));
    Odrv4 I__10387 (
            .O(N__47462),
            .I(\current_shift_inst.control_input_axb_19 ));
    InMux I__10386 (
            .O(N__47459),
            .I(N__47456));
    LocalMux I__10385 (
            .O(N__47456),
            .I(N__47453));
    Span4Mux_v I__10384 (
            .O(N__47453),
            .I(N__47450));
    Odrv4 I__10383 (
            .O(N__47450),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__10382 (
            .O(N__47447),
            .I(\current_shift_inst.control_input_cry_18 ));
    InMux I__10381 (
            .O(N__47444),
            .I(N__47441));
    LocalMux I__10380 (
            .O(N__47441),
            .I(\current_shift_inst.control_input_axb_20 ));
    InMux I__10379 (
            .O(N__47438),
            .I(N__47435));
    LocalMux I__10378 (
            .O(N__47435),
            .I(N__47432));
    Span4Mux_v I__10377 (
            .O(N__47432),
            .I(N__47429));
    Odrv4 I__10376 (
            .O(N__47429),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__10375 (
            .O(N__47426),
            .I(\current_shift_inst.control_input_cry_19 ));
    InMux I__10374 (
            .O(N__47423),
            .I(N__47420));
    LocalMux I__10373 (
            .O(N__47420),
            .I(\current_shift_inst.control_input_axb_21 ));
    InMux I__10372 (
            .O(N__47417),
            .I(N__47414));
    LocalMux I__10371 (
            .O(N__47414),
            .I(N__47411));
    Span4Mux_h I__10370 (
            .O(N__47411),
            .I(N__47408));
    Odrv4 I__10369 (
            .O(N__47408),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__10368 (
            .O(N__47405),
            .I(\current_shift_inst.control_input_cry_20 ));
    InMux I__10367 (
            .O(N__47402),
            .I(N__47399));
    LocalMux I__10366 (
            .O(N__47399),
            .I(N__47396));
    Odrv4 I__10365 (
            .O(N__47396),
            .I(\current_shift_inst.control_input_axb_22 ));
    InMux I__10364 (
            .O(N__47393),
            .I(N__47390));
    LocalMux I__10363 (
            .O(N__47390),
            .I(N__47387));
    Span4Mux_h I__10362 (
            .O(N__47387),
            .I(N__47384));
    Odrv4 I__10361 (
            .O(N__47384),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__10360 (
            .O(N__47381),
            .I(\current_shift_inst.control_input_cry_21 ));
    InMux I__10359 (
            .O(N__47378),
            .I(N__47375));
    LocalMux I__10358 (
            .O(N__47375),
            .I(\current_shift_inst.control_input_axb_23 ));
    InMux I__10357 (
            .O(N__47372),
            .I(N__47369));
    LocalMux I__10356 (
            .O(N__47369),
            .I(N__47366));
    Span4Mux_h I__10355 (
            .O(N__47366),
            .I(N__47363));
    Odrv4 I__10354 (
            .O(N__47363),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__10353 (
            .O(N__47360),
            .I(\current_shift_inst.control_input_cry_22 ));
    InMux I__10352 (
            .O(N__47357),
            .I(N__47354));
    LocalMux I__10351 (
            .O(N__47354),
            .I(N__47351));
    Span4Mux_v I__10350 (
            .O(N__47351),
            .I(N__47348));
    Odrv4 I__10349 (
            .O(N__47348),
            .I(\current_shift_inst.control_input_axb_24 ));
    InMux I__10348 (
            .O(N__47345),
            .I(N__47342));
    LocalMux I__10347 (
            .O(N__47342),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__10346 (
            .O(N__47339),
            .I(N__47336));
    LocalMux I__10345 (
            .O(N__47336),
            .I(N__47333));
    Span4Mux_h I__10344 (
            .O(N__47333),
            .I(N__47330));
    Odrv4 I__10343 (
            .O(N__47330),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__10342 (
            .O(N__47327),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__10341 (
            .O(N__47324),
            .I(N__47321));
    LocalMux I__10340 (
            .O(N__47321),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__10339 (
            .O(N__47318),
            .I(N__47315));
    LocalMux I__10338 (
            .O(N__47315),
            .I(N__47312));
    Span4Mux_v I__10337 (
            .O(N__47312),
            .I(N__47309));
    Odrv4 I__10336 (
            .O(N__47309),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__10335 (
            .O(N__47306),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__10334 (
            .O(N__47303),
            .I(N__47300));
    LocalMux I__10333 (
            .O(N__47300),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__10332 (
            .O(N__47297),
            .I(N__47294));
    LocalMux I__10331 (
            .O(N__47294),
            .I(N__47291));
    Span4Mux_v I__10330 (
            .O(N__47291),
            .I(N__47288));
    Odrv4 I__10329 (
            .O(N__47288),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__10328 (
            .O(N__47285),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__10327 (
            .O(N__47282),
            .I(N__47279));
    LocalMux I__10326 (
            .O(N__47279),
            .I(N__47276));
    Odrv4 I__10325 (
            .O(N__47276),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__10324 (
            .O(N__47273),
            .I(N__47270));
    LocalMux I__10323 (
            .O(N__47270),
            .I(N__47267));
    Span4Mux_h I__10322 (
            .O(N__47267),
            .I(N__47264));
    Odrv4 I__10321 (
            .O(N__47264),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__10320 (
            .O(N__47261),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__10319 (
            .O(N__47258),
            .I(N__47255));
    LocalMux I__10318 (
            .O(N__47255),
            .I(N__47252));
    Odrv4 I__10317 (
            .O(N__47252),
            .I(\current_shift_inst.control_input_axb_13 ));
    InMux I__10316 (
            .O(N__47249),
            .I(N__47246));
    LocalMux I__10315 (
            .O(N__47246),
            .I(N__47243));
    Span4Mux_h I__10314 (
            .O(N__47243),
            .I(N__47240));
    Odrv4 I__10313 (
            .O(N__47240),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__10312 (
            .O(N__47237),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__10311 (
            .O(N__47234),
            .I(N__47231));
    LocalMux I__10310 (
            .O(N__47231),
            .I(N__47228));
    Odrv4 I__10309 (
            .O(N__47228),
            .I(\current_shift_inst.control_input_axb_14 ));
    InMux I__10308 (
            .O(N__47225),
            .I(N__47222));
    LocalMux I__10307 (
            .O(N__47222),
            .I(N__47219));
    Span4Mux_h I__10306 (
            .O(N__47219),
            .I(N__47216));
    Odrv4 I__10305 (
            .O(N__47216),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__10304 (
            .O(N__47213),
            .I(\current_shift_inst.control_input_cry_13 ));
    InMux I__10303 (
            .O(N__47210),
            .I(N__47207));
    LocalMux I__10302 (
            .O(N__47207),
            .I(\current_shift_inst.control_input_axb_15 ));
    InMux I__10301 (
            .O(N__47204),
            .I(N__47201));
    LocalMux I__10300 (
            .O(N__47201),
            .I(N__47198));
    Span4Mux_h I__10299 (
            .O(N__47198),
            .I(N__47195));
    Odrv4 I__10298 (
            .O(N__47195),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__10297 (
            .O(N__47192),
            .I(\current_shift_inst.control_input_cry_14 ));
    InMux I__10296 (
            .O(N__47189),
            .I(N__47186));
    LocalMux I__10295 (
            .O(N__47186),
            .I(N__47183));
    Odrv4 I__10294 (
            .O(N__47183),
            .I(\current_shift_inst.control_input_axb_16 ));
    InMux I__10293 (
            .O(N__47180),
            .I(N__47177));
    LocalMux I__10292 (
            .O(N__47177),
            .I(N__47174));
    Span4Mux_h I__10291 (
            .O(N__47174),
            .I(N__47171));
    Odrv4 I__10290 (
            .O(N__47171),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__10289 (
            .O(N__47168),
            .I(bfn_17_21_0_));
    InMux I__10288 (
            .O(N__47165),
            .I(N__47162));
    LocalMux I__10287 (
            .O(N__47162),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__10286 (
            .O(N__47159),
            .I(N__47156));
    LocalMux I__10285 (
            .O(N__47156),
            .I(N__47153));
    Span4Mux_h I__10284 (
            .O(N__47153),
            .I(N__47150));
    Odrv4 I__10283 (
            .O(N__47150),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__10282 (
            .O(N__47147),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__10281 (
            .O(N__47144),
            .I(N__47141));
    LocalMux I__10280 (
            .O(N__47141),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__10279 (
            .O(N__47138),
            .I(N__47135));
    LocalMux I__10278 (
            .O(N__47135),
            .I(N__47132));
    Span4Mux_v I__10277 (
            .O(N__47132),
            .I(N__47129));
    Odrv4 I__10276 (
            .O(N__47129),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__10275 (
            .O(N__47126),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__10274 (
            .O(N__47123),
            .I(N__47120));
    LocalMux I__10273 (
            .O(N__47120),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__10272 (
            .O(N__47117),
            .I(N__47114));
    LocalMux I__10271 (
            .O(N__47114),
            .I(N__47111));
    Span4Mux_v I__10270 (
            .O(N__47111),
            .I(N__47108));
    Odrv4 I__10269 (
            .O(N__47108),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__10268 (
            .O(N__47105),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__10267 (
            .O(N__47102),
            .I(N__47099));
    LocalMux I__10266 (
            .O(N__47099),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__10265 (
            .O(N__47096),
            .I(N__47093));
    LocalMux I__10264 (
            .O(N__47093),
            .I(N__47090));
    Span4Mux_h I__10263 (
            .O(N__47090),
            .I(N__47087));
    Odrv4 I__10262 (
            .O(N__47087),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__10261 (
            .O(N__47084),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__10260 (
            .O(N__47081),
            .I(N__47078));
    LocalMux I__10259 (
            .O(N__47078),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__10258 (
            .O(N__47075),
            .I(N__47072));
    LocalMux I__10257 (
            .O(N__47072),
            .I(N__47069));
    Span4Mux_h I__10256 (
            .O(N__47069),
            .I(N__47066));
    Odrv4 I__10255 (
            .O(N__47066),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__10254 (
            .O(N__47063),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__10253 (
            .O(N__47060),
            .I(N__47057));
    LocalMux I__10252 (
            .O(N__47057),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__10251 (
            .O(N__47054),
            .I(N__47051));
    LocalMux I__10250 (
            .O(N__47051),
            .I(N__47048));
    Span4Mux_h I__10249 (
            .O(N__47048),
            .I(N__47045));
    Odrv4 I__10248 (
            .O(N__47045),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__10247 (
            .O(N__47042),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__10246 (
            .O(N__47039),
            .I(N__47036));
    LocalMux I__10245 (
            .O(N__47036),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__10244 (
            .O(N__47033),
            .I(N__47030));
    LocalMux I__10243 (
            .O(N__47030),
            .I(N__47027));
    Span4Mux_h I__10242 (
            .O(N__47027),
            .I(N__47024));
    Odrv4 I__10241 (
            .O(N__47024),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__10240 (
            .O(N__47021),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__10239 (
            .O(N__47018),
            .I(N__47015));
    LocalMux I__10238 (
            .O(N__47015),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__10237 (
            .O(N__47012),
            .I(N__47009));
    LocalMux I__10236 (
            .O(N__47009),
            .I(N__47006));
    Span4Mux_h I__10235 (
            .O(N__47006),
            .I(N__47003));
    Odrv4 I__10234 (
            .O(N__47003),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__10233 (
            .O(N__47000),
            .I(bfn_17_20_0_));
    InMux I__10232 (
            .O(N__46997),
            .I(N__46994));
    LocalMux I__10231 (
            .O(N__46994),
            .I(N__46991));
    Span12Mux_h I__10230 (
            .O(N__46991),
            .I(N__46988));
    Odrv12 I__10229 (
            .O(N__46988),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__10228 (
            .O(N__46985),
            .I(N__46982));
    LocalMux I__10227 (
            .O(N__46982),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__10226 (
            .O(N__46979),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    CascadeMux I__10225 (
            .O(N__46976),
            .I(N__46973));
    InMux I__10224 (
            .O(N__46973),
            .I(N__46970));
    LocalMux I__10223 (
            .O(N__46970),
            .I(N__46967));
    Odrv12 I__10222 (
            .O(N__46967),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__10221 (
            .O(N__46964),
            .I(N__46961));
    LocalMux I__10220 (
            .O(N__46961),
            .I(N__46958));
    Span4Mux_h I__10219 (
            .O(N__46958),
            .I(N__46955));
    Odrv4 I__10218 (
            .O(N__46955),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__10217 (
            .O(N__46952),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__10216 (
            .O(N__46949),
            .I(N__46946));
    LocalMux I__10215 (
            .O(N__46946),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__10214 (
            .O(N__46943),
            .I(N__46940));
    LocalMux I__10213 (
            .O(N__46940),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__10212 (
            .O(N__46937),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    CascadeMux I__10211 (
            .O(N__46934),
            .I(N__46931));
    InMux I__10210 (
            .O(N__46931),
            .I(N__46928));
    LocalMux I__10209 (
            .O(N__46928),
            .I(N__46925));
    Span4Mux_v I__10208 (
            .O(N__46925),
            .I(N__46922));
    Odrv4 I__10207 (
            .O(N__46922),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__10206 (
            .O(N__46919),
            .I(N__46916));
    LocalMux I__10205 (
            .O(N__46916),
            .I(N__46913));
    Odrv4 I__10204 (
            .O(N__46913),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__10203 (
            .O(N__46910),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__10202 (
            .O(N__46907),
            .I(N__46904));
    LocalMux I__10201 (
            .O(N__46904),
            .I(N__46901));
    Odrv12 I__10200 (
            .O(N__46901),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__10199 (
            .O(N__46898),
            .I(N__46895));
    LocalMux I__10198 (
            .O(N__46895),
            .I(N__46892));
    Sp12to4 I__10197 (
            .O(N__46892),
            .I(N__46889));
    Odrv12 I__10196 (
            .O(N__46889),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__10195 (
            .O(N__46886),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    CascadeMux I__10194 (
            .O(N__46883),
            .I(N__46880));
    InMux I__10193 (
            .O(N__46880),
            .I(N__46877));
    LocalMux I__10192 (
            .O(N__46877),
            .I(N__46874));
    Span4Mux_h I__10191 (
            .O(N__46874),
            .I(N__46871));
    Odrv4 I__10190 (
            .O(N__46871),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__10189 (
            .O(N__46868),
            .I(N__46865));
    LocalMux I__10188 (
            .O(N__46865),
            .I(N__46862));
    Odrv4 I__10187 (
            .O(N__46862),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__10186 (
            .O(N__46859),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__10185 (
            .O(N__46856),
            .I(N__46853));
    LocalMux I__10184 (
            .O(N__46853),
            .I(N__46850));
    Span4Mux_h I__10183 (
            .O(N__46850),
            .I(N__46847));
    Odrv4 I__10182 (
            .O(N__46847),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__10181 (
            .O(N__46844),
            .I(N__46841));
    LocalMux I__10180 (
            .O(N__46841),
            .I(N__46838));
    Odrv4 I__10179 (
            .O(N__46838),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__10178 (
            .O(N__46835),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__10177 (
            .O(N__46832),
            .I(N__46829));
    LocalMux I__10176 (
            .O(N__46829),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__10175 (
            .O(N__46826),
            .I(N__46821));
    InMux I__10174 (
            .O(N__46825),
            .I(N__46818));
    InMux I__10173 (
            .O(N__46824),
            .I(N__46815));
    InMux I__10172 (
            .O(N__46821),
            .I(N__46812));
    LocalMux I__10171 (
            .O(N__46818),
            .I(\current_shift_inst.N_1619_i ));
    LocalMux I__10170 (
            .O(N__46815),
            .I(\current_shift_inst.N_1619_i ));
    LocalMux I__10169 (
            .O(N__46812),
            .I(\current_shift_inst.N_1619_i ));
    InMux I__10168 (
            .O(N__46805),
            .I(N__46802));
    LocalMux I__10167 (
            .O(N__46802),
            .I(N__46799));
    Span4Mux_h I__10166 (
            .O(N__46799),
            .I(N__46796));
    Odrv4 I__10165 (
            .O(N__46796),
            .I(\current_shift_inst.control_input_1 ));
    InMux I__10164 (
            .O(N__46793),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    CascadeMux I__10163 (
            .O(N__46790),
            .I(N__46787));
    InMux I__10162 (
            .O(N__46787),
            .I(N__46784));
    LocalMux I__10161 (
            .O(N__46784),
            .I(N__46781));
    Span4Mux_h I__10160 (
            .O(N__46781),
            .I(N__46778));
    Odrv4 I__10159 (
            .O(N__46778),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    InMux I__10158 (
            .O(N__46775),
            .I(N__46772));
    LocalMux I__10157 (
            .O(N__46772),
            .I(N__46769));
    Span4Mux_v I__10156 (
            .O(N__46769),
            .I(N__46766));
    Odrv4 I__10155 (
            .O(N__46766),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__10154 (
            .O(N__46763),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__10153 (
            .O(N__46760),
            .I(N__46757));
    LocalMux I__10152 (
            .O(N__46757),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__10151 (
            .O(N__46754),
            .I(N__46751));
    LocalMux I__10150 (
            .O(N__46751),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__10149 (
            .O(N__46748),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    CascadeMux I__10148 (
            .O(N__46745),
            .I(N__46742));
    InMux I__10147 (
            .O(N__46742),
            .I(N__46739));
    LocalMux I__10146 (
            .O(N__46739),
            .I(N__46736));
    Odrv12 I__10145 (
            .O(N__46736),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__10144 (
            .O(N__46733),
            .I(N__46730));
    LocalMux I__10143 (
            .O(N__46730),
            .I(N__46727));
    Span4Mux_h I__10142 (
            .O(N__46727),
            .I(N__46724));
    Span4Mux_v I__10141 (
            .O(N__46724),
            .I(N__46721));
    Odrv4 I__10140 (
            .O(N__46721),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__10139 (
            .O(N__46718),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__10138 (
            .O(N__46715),
            .I(N__46712));
    LocalMux I__10137 (
            .O(N__46712),
            .I(N__46709));
    Odrv4 I__10136 (
            .O(N__46709),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__10135 (
            .O(N__46706),
            .I(N__46703));
    LocalMux I__10134 (
            .O(N__46703),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__10133 (
            .O(N__46700),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    CascadeMux I__10132 (
            .O(N__46697),
            .I(N__46694));
    InMux I__10131 (
            .O(N__46694),
            .I(N__46691));
    LocalMux I__10130 (
            .O(N__46691),
            .I(N__46688));
    Span4Mux_h I__10129 (
            .O(N__46688),
            .I(N__46685));
    Odrv4 I__10128 (
            .O(N__46685),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__10127 (
            .O(N__46682),
            .I(N__46679));
    LocalMux I__10126 (
            .O(N__46679),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__10125 (
            .O(N__46676),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__10124 (
            .O(N__46673),
            .I(N__46670));
    LocalMux I__10123 (
            .O(N__46670),
            .I(N__46667));
    Span4Mux_h I__10122 (
            .O(N__46667),
            .I(N__46664));
    Odrv4 I__10121 (
            .O(N__46664),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__10120 (
            .O(N__46661),
            .I(N__46658));
    LocalMux I__10119 (
            .O(N__46658),
            .I(N__46655));
    Span4Mux_v I__10118 (
            .O(N__46655),
            .I(N__46652));
    Odrv4 I__10117 (
            .O(N__46652),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__10116 (
            .O(N__46649),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    CascadeMux I__10115 (
            .O(N__46646),
            .I(N__46643));
    InMux I__10114 (
            .O(N__46643),
            .I(N__46640));
    LocalMux I__10113 (
            .O(N__46640),
            .I(N__46637));
    Odrv4 I__10112 (
            .O(N__46637),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__10111 (
            .O(N__46634),
            .I(N__46631));
    LocalMux I__10110 (
            .O(N__46631),
            .I(N__46628));
    Span4Mux_v I__10109 (
            .O(N__46628),
            .I(N__46625));
    Odrv4 I__10108 (
            .O(N__46625),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__10107 (
            .O(N__46622),
            .I(bfn_17_18_0_));
    CascadeMux I__10106 (
            .O(N__46619),
            .I(N__46616));
    InMux I__10105 (
            .O(N__46616),
            .I(N__46613));
    LocalMux I__10104 (
            .O(N__46613),
            .I(N__46610));
    Span4Mux_h I__10103 (
            .O(N__46610),
            .I(N__46607));
    Odrv4 I__10102 (
            .O(N__46607),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    InMux I__10101 (
            .O(N__46604),
            .I(N__46601));
    LocalMux I__10100 (
            .O(N__46601),
            .I(N__46598));
    Odrv4 I__10099 (
            .O(N__46598),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__10098 (
            .O(N__46595),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__10097 (
            .O(N__46592),
            .I(N__46589));
    LocalMux I__10096 (
            .O(N__46589),
            .I(N__46586));
    Odrv12 I__10095 (
            .O(N__46586),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    InMux I__10094 (
            .O(N__46583),
            .I(N__46580));
    LocalMux I__10093 (
            .O(N__46580),
            .I(N__46577));
    Span4Mux_v I__10092 (
            .O(N__46577),
            .I(N__46574));
    Odrv4 I__10091 (
            .O(N__46574),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__10090 (
            .O(N__46571),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    CascadeMux I__10089 (
            .O(N__46568),
            .I(N__46565));
    InMux I__10088 (
            .O(N__46565),
            .I(N__46562));
    LocalMux I__10087 (
            .O(N__46562),
            .I(N__46559));
    Odrv4 I__10086 (
            .O(N__46559),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    InMux I__10085 (
            .O(N__46556),
            .I(N__46553));
    LocalMux I__10084 (
            .O(N__46553),
            .I(N__46550));
    Span4Mux_v I__10083 (
            .O(N__46550),
            .I(N__46547));
    Odrv4 I__10082 (
            .O(N__46547),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__10081 (
            .O(N__46544),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__10080 (
            .O(N__46541),
            .I(N__46538));
    LocalMux I__10079 (
            .O(N__46538),
            .I(N__46535));
    Span4Mux_h I__10078 (
            .O(N__46535),
            .I(N__46532));
    Odrv4 I__10077 (
            .O(N__46532),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    InMux I__10076 (
            .O(N__46529),
            .I(N__46526));
    LocalMux I__10075 (
            .O(N__46526),
            .I(N__46523));
    Span4Mux_v I__10074 (
            .O(N__46523),
            .I(N__46520));
    Odrv4 I__10073 (
            .O(N__46520),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__10072 (
            .O(N__46517),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    CascadeMux I__10071 (
            .O(N__46514),
            .I(N__46511));
    InMux I__10070 (
            .O(N__46511),
            .I(N__46508));
    LocalMux I__10069 (
            .O(N__46508),
            .I(N__46505));
    Odrv4 I__10068 (
            .O(N__46505),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__10067 (
            .O(N__46502),
            .I(N__46499));
    LocalMux I__10066 (
            .O(N__46499),
            .I(N__46496));
    Span4Mux_v I__10065 (
            .O(N__46496),
            .I(N__46493));
    Odrv4 I__10064 (
            .O(N__46493),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__10063 (
            .O(N__46490),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__10062 (
            .O(N__46487),
            .I(N__46484));
    LocalMux I__10061 (
            .O(N__46484),
            .I(N__46481));
    Odrv12 I__10060 (
            .O(N__46481),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__10059 (
            .O(N__46478),
            .I(N__46475));
    LocalMux I__10058 (
            .O(N__46475),
            .I(N__46472));
    Odrv4 I__10057 (
            .O(N__46472),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__10056 (
            .O(N__46469),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    CascadeMux I__10055 (
            .O(N__46466),
            .I(N__46463));
    InMux I__10054 (
            .O(N__46463),
            .I(N__46460));
    LocalMux I__10053 (
            .O(N__46460),
            .I(N__46457));
    Span4Mux_h I__10052 (
            .O(N__46457),
            .I(N__46454));
    Span4Mux_h I__10051 (
            .O(N__46454),
            .I(N__46451));
    Odrv4 I__10050 (
            .O(N__46451),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__10049 (
            .O(N__46448),
            .I(N__46445));
    LocalMux I__10048 (
            .O(N__46445),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__10047 (
            .O(N__46442),
            .I(bfn_17_17_0_));
    InMux I__10046 (
            .O(N__46439),
            .I(N__46436));
    LocalMux I__10045 (
            .O(N__46436),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__10044 (
            .O(N__46433),
            .I(N__46430));
    LocalMux I__10043 (
            .O(N__46430),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    CascadeMux I__10042 (
            .O(N__46427),
            .I(N__46422));
    InMux I__10041 (
            .O(N__46426),
            .I(N__46414));
    InMux I__10040 (
            .O(N__46425),
            .I(N__46414));
    InMux I__10039 (
            .O(N__46422),
            .I(N__46409));
    InMux I__10038 (
            .O(N__46421),
            .I(N__46409));
    InMux I__10037 (
            .O(N__46420),
            .I(N__46406));
    CascadeMux I__10036 (
            .O(N__46419),
            .I(N__46403));
    LocalMux I__10035 (
            .O(N__46414),
            .I(N__46400));
    LocalMux I__10034 (
            .O(N__46409),
            .I(N__46397));
    LocalMux I__10033 (
            .O(N__46406),
            .I(N__46394));
    InMux I__10032 (
            .O(N__46403),
            .I(N__46391));
    Span4Mux_h I__10031 (
            .O(N__46400),
            .I(N__46388));
    Span4Mux_h I__10030 (
            .O(N__46397),
            .I(N__46381));
    Span4Mux_h I__10029 (
            .O(N__46394),
            .I(N__46381));
    LocalMux I__10028 (
            .O(N__46391),
            .I(N__46381));
    Odrv4 I__10027 (
            .O(N__46388),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__10026 (
            .O(N__46381),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__10025 (
            .O(N__46376),
            .I(N__46373));
    InMux I__10024 (
            .O(N__46373),
            .I(N__46370));
    LocalMux I__10023 (
            .O(N__46370),
            .I(N__46367));
    Span4Mux_v I__10022 (
            .O(N__46367),
            .I(N__46364));
    Span4Mux_h I__10021 (
            .O(N__46364),
            .I(N__46361));
    Odrv4 I__10020 (
            .O(N__46361),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__10019 (
            .O(N__46358),
            .I(N__46355));
    LocalMux I__10018 (
            .O(N__46355),
            .I(N__46352));
    Span4Mux_v I__10017 (
            .O(N__46352),
            .I(N__46349));
    Odrv4 I__10016 (
            .O(N__46349),
            .I(\current_shift_inst.un38_control_input_0_s0_3 ));
    InMux I__10015 (
            .O(N__46346),
            .I(\current_shift_inst.un38_control_input_cry_2_s0 ));
    CascadeMux I__10014 (
            .O(N__46343),
            .I(N__46340));
    InMux I__10013 (
            .O(N__46340),
            .I(N__46337));
    LocalMux I__10012 (
            .O(N__46337),
            .I(N__46334));
    Span4Mux_h I__10011 (
            .O(N__46334),
            .I(N__46331));
    Odrv4 I__10010 (
            .O(N__46331),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ));
    InMux I__10009 (
            .O(N__46328),
            .I(N__46325));
    LocalMux I__10008 (
            .O(N__46325),
            .I(N__46322));
    Span4Mux_v I__10007 (
            .O(N__46322),
            .I(N__46319));
    Odrv4 I__10006 (
            .O(N__46319),
            .I(\current_shift_inst.un38_control_input_0_s0_4 ));
    InMux I__10005 (
            .O(N__46316),
            .I(\current_shift_inst.un38_control_input_cry_3_s0 ));
    InMux I__10004 (
            .O(N__46313),
            .I(N__46310));
    LocalMux I__10003 (
            .O(N__46310),
            .I(N__46307));
    Span4Mux_v I__10002 (
            .O(N__46307),
            .I(N__46304));
    Odrv4 I__10001 (
            .O(N__46304),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ));
    InMux I__10000 (
            .O(N__46301),
            .I(N__46298));
    LocalMux I__9999 (
            .O(N__46298),
            .I(N__46295));
    Sp12to4 I__9998 (
            .O(N__46295),
            .I(N__46292));
    Odrv12 I__9997 (
            .O(N__46292),
            .I(\current_shift_inst.un38_control_input_0_s0_5 ));
    InMux I__9996 (
            .O(N__46289),
            .I(\current_shift_inst.un38_control_input_cry_4_s0 ));
    CascadeMux I__9995 (
            .O(N__46286),
            .I(N__46283));
    InMux I__9994 (
            .O(N__46283),
            .I(N__46280));
    LocalMux I__9993 (
            .O(N__46280),
            .I(N__46277));
    Span4Mux_h I__9992 (
            .O(N__46277),
            .I(N__46274));
    Odrv4 I__9991 (
            .O(N__46274),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    InMux I__9990 (
            .O(N__46271),
            .I(N__46268));
    LocalMux I__9989 (
            .O(N__46268),
            .I(N__46265));
    Span4Mux_v I__9988 (
            .O(N__46265),
            .I(N__46262));
    Odrv4 I__9987 (
            .O(N__46262),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__9986 (
            .O(N__46259),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__9985 (
            .O(N__46256),
            .I(N__46253));
    LocalMux I__9984 (
            .O(N__46253),
            .I(N__46250));
    Span4Mux_v I__9983 (
            .O(N__46250),
            .I(N__46247));
    Odrv4 I__9982 (
            .O(N__46247),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    InMux I__9981 (
            .O(N__46244),
            .I(N__46241));
    LocalMux I__9980 (
            .O(N__46241),
            .I(N__46238));
    Span4Mux_v I__9979 (
            .O(N__46238),
            .I(N__46235));
    Odrv4 I__9978 (
            .O(N__46235),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__9977 (
            .O(N__46232),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    CascadeMux I__9976 (
            .O(N__46229),
            .I(N__46226));
    InMux I__9975 (
            .O(N__46226),
            .I(N__46223));
    LocalMux I__9974 (
            .O(N__46223),
            .I(N__46220));
    Span4Mux_h I__9973 (
            .O(N__46220),
            .I(N__46217));
    Span4Mux_v I__9972 (
            .O(N__46217),
            .I(N__46214));
    Odrv4 I__9971 (
            .O(N__46214),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    InMux I__9970 (
            .O(N__46211),
            .I(N__46208));
    LocalMux I__9969 (
            .O(N__46208),
            .I(N__46205));
    Span4Mux_v I__9968 (
            .O(N__46205),
            .I(N__46202));
    Odrv4 I__9967 (
            .O(N__46202),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__9966 (
            .O(N__46199),
            .I(bfn_17_16_0_));
    InMux I__9965 (
            .O(N__46196),
            .I(N__46193));
    LocalMux I__9964 (
            .O(N__46193),
            .I(N__46190));
    Span4Mux_v I__9963 (
            .O(N__46190),
            .I(N__46187));
    Odrv4 I__9962 (
            .O(N__46187),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    InMux I__9961 (
            .O(N__46184),
            .I(N__46181));
    LocalMux I__9960 (
            .O(N__46181),
            .I(N__46178));
    Span4Mux_v I__9959 (
            .O(N__46178),
            .I(N__46175));
    Odrv4 I__9958 (
            .O(N__46175),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__9957 (
            .O(N__46172),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    CascadeMux I__9956 (
            .O(N__46169),
            .I(N__46166));
    InMux I__9955 (
            .O(N__46166),
            .I(N__46162));
    InMux I__9954 (
            .O(N__46165),
            .I(N__46159));
    LocalMux I__9953 (
            .O(N__46162),
            .I(N__46155));
    LocalMux I__9952 (
            .O(N__46159),
            .I(N__46152));
    InMux I__9951 (
            .O(N__46158),
            .I(N__46149));
    Span4Mux_v I__9950 (
            .O(N__46155),
            .I(N__46146));
    Span4Mux_h I__9949 (
            .O(N__46152),
            .I(N__46143));
    LocalMux I__9948 (
            .O(N__46149),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__9947 (
            .O(N__46146),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__9946 (
            .O(N__46143),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__9945 (
            .O(N__46136),
            .I(bfn_17_14_0_));
    CascadeMux I__9944 (
            .O(N__46133),
            .I(N__46129));
    CascadeMux I__9943 (
            .O(N__46132),
            .I(N__46126));
    InMux I__9942 (
            .O(N__46129),
            .I(N__46122));
    InMux I__9941 (
            .O(N__46126),
            .I(N__46119));
    InMux I__9940 (
            .O(N__46125),
            .I(N__46116));
    LocalMux I__9939 (
            .O(N__46122),
            .I(N__46113));
    LocalMux I__9938 (
            .O(N__46119),
            .I(N__46110));
    LocalMux I__9937 (
            .O(N__46116),
            .I(N__46105));
    Span4Mux_v I__9936 (
            .O(N__46113),
            .I(N__46105));
    Span4Mux_h I__9935 (
            .O(N__46110),
            .I(N__46102));
    Odrv4 I__9934 (
            .O(N__46105),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__9933 (
            .O(N__46102),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__9932 (
            .O(N__46097),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__9931 (
            .O(N__46094),
            .I(N__46088));
    InMux I__9930 (
            .O(N__46093),
            .I(N__46088));
    LocalMux I__9929 (
            .O(N__46088),
            .I(N__46084));
    InMux I__9928 (
            .O(N__46087),
            .I(N__46081));
    Span4Mux_h I__9927 (
            .O(N__46084),
            .I(N__46078));
    LocalMux I__9926 (
            .O(N__46081),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__9925 (
            .O(N__46078),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__9924 (
            .O(N__46073),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__9923 (
            .O(N__46070),
            .I(N__46064));
    InMux I__9922 (
            .O(N__46069),
            .I(N__46064));
    LocalMux I__9921 (
            .O(N__46064),
            .I(N__46060));
    InMux I__9920 (
            .O(N__46063),
            .I(N__46057));
    Span4Mux_h I__9919 (
            .O(N__46060),
            .I(N__46054));
    LocalMux I__9918 (
            .O(N__46057),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__9917 (
            .O(N__46054),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__9916 (
            .O(N__46049),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    CascadeMux I__9915 (
            .O(N__46046),
            .I(N__46043));
    InMux I__9914 (
            .O(N__46043),
            .I(N__46040));
    LocalMux I__9913 (
            .O(N__46040),
            .I(N__46037));
    Span4Mux_h I__9912 (
            .O(N__46037),
            .I(N__46033));
    InMux I__9911 (
            .O(N__46036),
            .I(N__46030));
    Span4Mux_h I__9910 (
            .O(N__46033),
            .I(N__46027));
    LocalMux I__9909 (
            .O(N__46030),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__9908 (
            .O(N__46027),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__9907 (
            .O(N__46022),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__9906 (
            .O(N__46019),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__9905 (
            .O(N__46016),
            .I(N__46013));
    InMux I__9904 (
            .O(N__46013),
            .I(N__46010));
    LocalMux I__9903 (
            .O(N__46010),
            .I(N__46006));
    InMux I__9902 (
            .O(N__46009),
            .I(N__46003));
    Span4Mux_h I__9901 (
            .O(N__46006),
            .I(N__46000));
    LocalMux I__9900 (
            .O(N__46003),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__9899 (
            .O(N__46000),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    InMux I__9898 (
            .O(N__45995),
            .I(N__45992));
    LocalMux I__9897 (
            .O(N__45992),
            .I(N__45989));
    Span4Mux_v I__9896 (
            .O(N__45989),
            .I(N__45986));
    Odrv4 I__9895 (
            .O(N__45986),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__9894 (
            .O(N__45983),
            .I(N__45980));
    InMux I__9893 (
            .O(N__45980),
            .I(N__45976));
    CascadeMux I__9892 (
            .O(N__45979),
            .I(N__45973));
    LocalMux I__9891 (
            .O(N__45976),
            .I(N__45970));
    InMux I__9890 (
            .O(N__45973),
            .I(N__45967));
    Span4Mux_v I__9889 (
            .O(N__45970),
            .I(N__45962));
    LocalMux I__9888 (
            .O(N__45967),
            .I(N__45962));
    Odrv4 I__9887 (
            .O(N__45962),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__9886 (
            .O(N__45959),
            .I(N__45956));
    InMux I__9885 (
            .O(N__45956),
            .I(N__45953));
    LocalMux I__9884 (
            .O(N__45953),
            .I(N__45950));
    Span4Mux_h I__9883 (
            .O(N__45950),
            .I(N__45947));
    Odrv4 I__9882 (
            .O(N__45947),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    CascadeMux I__9881 (
            .O(N__45944),
            .I(N__45940));
    InMux I__9880 (
            .O(N__45943),
            .I(N__45935));
    InMux I__9879 (
            .O(N__45940),
            .I(N__45935));
    LocalMux I__9878 (
            .O(N__45935),
            .I(N__45932));
    Span4Mux_v I__9877 (
            .O(N__45932),
            .I(N__45927));
    InMux I__9876 (
            .O(N__45931),
            .I(N__45924));
    InMux I__9875 (
            .O(N__45930),
            .I(N__45921));
    Span4Mux_h I__9874 (
            .O(N__45927),
            .I(N__45916));
    LocalMux I__9873 (
            .O(N__45924),
            .I(N__45916));
    LocalMux I__9872 (
            .O(N__45921),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__9871 (
            .O(N__45916),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    InMux I__9870 (
            .O(N__45911),
            .I(N__45905));
    InMux I__9869 (
            .O(N__45910),
            .I(N__45905));
    LocalMux I__9868 (
            .O(N__45905),
            .I(N__45901));
    InMux I__9867 (
            .O(N__45904),
            .I(N__45898));
    Span4Mux_h I__9866 (
            .O(N__45901),
            .I(N__45895));
    LocalMux I__9865 (
            .O(N__45898),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__9864 (
            .O(N__45895),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__9863 (
            .O(N__45890),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__9862 (
            .O(N__45887),
            .I(N__45884));
    InMux I__9861 (
            .O(N__45884),
            .I(N__45879));
    InMux I__9860 (
            .O(N__45883),
            .I(N__45876));
    InMux I__9859 (
            .O(N__45882),
            .I(N__45873));
    LocalMux I__9858 (
            .O(N__45879),
            .I(N__45870));
    LocalMux I__9857 (
            .O(N__45876),
            .I(N__45867));
    LocalMux I__9856 (
            .O(N__45873),
            .I(N__45862));
    Span4Mux_v I__9855 (
            .O(N__45870),
            .I(N__45862));
    Span4Mux_h I__9854 (
            .O(N__45867),
            .I(N__45859));
    Odrv4 I__9853 (
            .O(N__45862),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__9852 (
            .O(N__45859),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__9851 (
            .O(N__45854),
            .I(bfn_17_13_0_));
    CascadeMux I__9850 (
            .O(N__45851),
            .I(N__45847));
    CascadeMux I__9849 (
            .O(N__45850),
            .I(N__45844));
    InMux I__9848 (
            .O(N__45847),
            .I(N__45840));
    InMux I__9847 (
            .O(N__45844),
            .I(N__45837));
    InMux I__9846 (
            .O(N__45843),
            .I(N__45834));
    LocalMux I__9845 (
            .O(N__45840),
            .I(N__45831));
    LocalMux I__9844 (
            .O(N__45837),
            .I(N__45828));
    LocalMux I__9843 (
            .O(N__45834),
            .I(N__45823));
    Span4Mux_v I__9842 (
            .O(N__45831),
            .I(N__45823));
    Span4Mux_h I__9841 (
            .O(N__45828),
            .I(N__45820));
    Odrv4 I__9840 (
            .O(N__45823),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__9839 (
            .O(N__45820),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__9838 (
            .O(N__45815),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    CascadeMux I__9837 (
            .O(N__45812),
            .I(N__45809));
    InMux I__9836 (
            .O(N__45809),
            .I(N__45805));
    InMux I__9835 (
            .O(N__45808),
            .I(N__45802));
    LocalMux I__9834 (
            .O(N__45805),
            .I(N__45796));
    LocalMux I__9833 (
            .O(N__45802),
            .I(N__45796));
    InMux I__9832 (
            .O(N__45801),
            .I(N__45793));
    Span4Mux_h I__9831 (
            .O(N__45796),
            .I(N__45790));
    LocalMux I__9830 (
            .O(N__45793),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__9829 (
            .O(N__45790),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__9828 (
            .O(N__45785),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__9827 (
            .O(N__45782),
            .I(N__45776));
    InMux I__9826 (
            .O(N__45781),
            .I(N__45776));
    LocalMux I__9825 (
            .O(N__45776),
            .I(N__45772));
    InMux I__9824 (
            .O(N__45775),
            .I(N__45769));
    Span4Mux_h I__9823 (
            .O(N__45772),
            .I(N__45766));
    LocalMux I__9822 (
            .O(N__45769),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__9821 (
            .O(N__45766),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__9820 (
            .O(N__45761),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__9819 (
            .O(N__45758),
            .I(N__45755));
    InMux I__9818 (
            .O(N__45755),
            .I(N__45751));
    InMux I__9817 (
            .O(N__45754),
            .I(N__45748));
    LocalMux I__9816 (
            .O(N__45751),
            .I(N__45742));
    LocalMux I__9815 (
            .O(N__45748),
            .I(N__45742));
    InMux I__9814 (
            .O(N__45747),
            .I(N__45739));
    Span4Mux_h I__9813 (
            .O(N__45742),
            .I(N__45736));
    LocalMux I__9812 (
            .O(N__45739),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__9811 (
            .O(N__45736),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__9810 (
            .O(N__45731),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__9809 (
            .O(N__45728),
            .I(N__45724));
    CascadeMux I__9808 (
            .O(N__45727),
            .I(N__45721));
    InMux I__9807 (
            .O(N__45724),
            .I(N__45716));
    InMux I__9806 (
            .O(N__45721),
            .I(N__45716));
    LocalMux I__9805 (
            .O(N__45716),
            .I(N__45712));
    InMux I__9804 (
            .O(N__45715),
            .I(N__45709));
    Span4Mux_v I__9803 (
            .O(N__45712),
            .I(N__45706));
    LocalMux I__9802 (
            .O(N__45709),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__9801 (
            .O(N__45706),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__9800 (
            .O(N__45701),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__9799 (
            .O(N__45698),
            .I(N__45695));
    InMux I__9798 (
            .O(N__45695),
            .I(N__45691));
    InMux I__9797 (
            .O(N__45694),
            .I(N__45688));
    LocalMux I__9796 (
            .O(N__45691),
            .I(N__45682));
    LocalMux I__9795 (
            .O(N__45688),
            .I(N__45682));
    InMux I__9794 (
            .O(N__45687),
            .I(N__45679));
    Span4Mux_v I__9793 (
            .O(N__45682),
            .I(N__45676));
    LocalMux I__9792 (
            .O(N__45679),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__9791 (
            .O(N__45676),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__9790 (
            .O(N__45671),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__9789 (
            .O(N__45668),
            .I(N__45662));
    InMux I__9788 (
            .O(N__45667),
            .I(N__45662));
    LocalMux I__9787 (
            .O(N__45662),
            .I(N__45658));
    InMux I__9786 (
            .O(N__45661),
            .I(N__45655));
    Span4Mux_h I__9785 (
            .O(N__45658),
            .I(N__45652));
    LocalMux I__9784 (
            .O(N__45655),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__9783 (
            .O(N__45652),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__9782 (
            .O(N__45647),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__9781 (
            .O(N__45644),
            .I(N__45638));
    InMux I__9780 (
            .O(N__45643),
            .I(N__45638));
    LocalMux I__9779 (
            .O(N__45638),
            .I(N__45634));
    InMux I__9778 (
            .O(N__45637),
            .I(N__45631));
    Span4Mux_h I__9777 (
            .O(N__45634),
            .I(N__45628));
    LocalMux I__9776 (
            .O(N__45631),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__9775 (
            .O(N__45628),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__9774 (
            .O(N__45623),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__9773 (
            .O(N__45620),
            .I(N__45617));
    InMux I__9772 (
            .O(N__45617),
            .I(N__45612));
    InMux I__9771 (
            .O(N__45616),
            .I(N__45609));
    InMux I__9770 (
            .O(N__45615),
            .I(N__45606));
    LocalMux I__9769 (
            .O(N__45612),
            .I(N__45603));
    LocalMux I__9768 (
            .O(N__45609),
            .I(N__45600));
    LocalMux I__9767 (
            .O(N__45606),
            .I(N__45595));
    Span4Mux_v I__9766 (
            .O(N__45603),
            .I(N__45595));
    Span4Mux_h I__9765 (
            .O(N__45600),
            .I(N__45592));
    Odrv4 I__9764 (
            .O(N__45595),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__9763 (
            .O(N__45592),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__9762 (
            .O(N__45587),
            .I(bfn_17_12_0_));
    CascadeMux I__9761 (
            .O(N__45584),
            .I(N__45580));
    CascadeMux I__9760 (
            .O(N__45583),
            .I(N__45577));
    InMux I__9759 (
            .O(N__45580),
            .I(N__45574));
    InMux I__9758 (
            .O(N__45577),
            .I(N__45571));
    LocalMux I__9757 (
            .O(N__45574),
            .I(N__45567));
    LocalMux I__9756 (
            .O(N__45571),
            .I(N__45564));
    InMux I__9755 (
            .O(N__45570),
            .I(N__45561));
    Span4Mux_v I__9754 (
            .O(N__45567),
            .I(N__45558));
    Span4Mux_h I__9753 (
            .O(N__45564),
            .I(N__45555));
    LocalMux I__9752 (
            .O(N__45561),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__9751 (
            .O(N__45558),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__9750 (
            .O(N__45555),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__9749 (
            .O(N__45548),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__9748 (
            .O(N__45545),
            .I(N__45542));
    InMux I__9747 (
            .O(N__45542),
            .I(N__45538));
    InMux I__9746 (
            .O(N__45541),
            .I(N__45535));
    LocalMux I__9745 (
            .O(N__45538),
            .I(N__45529));
    LocalMux I__9744 (
            .O(N__45535),
            .I(N__45529));
    InMux I__9743 (
            .O(N__45534),
            .I(N__45526));
    Span4Mux_h I__9742 (
            .O(N__45529),
            .I(N__45523));
    LocalMux I__9741 (
            .O(N__45526),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__9740 (
            .O(N__45523),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__9739 (
            .O(N__45518),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__9738 (
            .O(N__45515),
            .I(N__45509));
    InMux I__9737 (
            .O(N__45514),
            .I(N__45509));
    LocalMux I__9736 (
            .O(N__45509),
            .I(N__45505));
    InMux I__9735 (
            .O(N__45508),
            .I(N__45502));
    Span4Mux_h I__9734 (
            .O(N__45505),
            .I(N__45499));
    LocalMux I__9733 (
            .O(N__45502),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__9732 (
            .O(N__45499),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__9731 (
            .O(N__45494),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__9730 (
            .O(N__45491),
            .I(N__45485));
    InMux I__9729 (
            .O(N__45490),
            .I(N__45485));
    LocalMux I__9728 (
            .O(N__45485),
            .I(N__45481));
    InMux I__9727 (
            .O(N__45484),
            .I(N__45478));
    Span4Mux_h I__9726 (
            .O(N__45481),
            .I(N__45475));
    LocalMux I__9725 (
            .O(N__45478),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__9724 (
            .O(N__45475),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__9723 (
            .O(N__45470),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__9722 (
            .O(N__45467),
            .I(N__45463));
    CascadeMux I__9721 (
            .O(N__45466),
            .I(N__45460));
    InMux I__9720 (
            .O(N__45463),
            .I(N__45455));
    InMux I__9719 (
            .O(N__45460),
            .I(N__45455));
    LocalMux I__9718 (
            .O(N__45455),
            .I(N__45451));
    InMux I__9717 (
            .O(N__45454),
            .I(N__45448));
    Span4Mux_h I__9716 (
            .O(N__45451),
            .I(N__45445));
    LocalMux I__9715 (
            .O(N__45448),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__9714 (
            .O(N__45445),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__9713 (
            .O(N__45440),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__9712 (
            .O(N__45437),
            .I(N__45433));
    CascadeMux I__9711 (
            .O(N__45436),
            .I(N__45430));
    InMux I__9710 (
            .O(N__45433),
            .I(N__45425));
    InMux I__9709 (
            .O(N__45430),
            .I(N__45425));
    LocalMux I__9708 (
            .O(N__45425),
            .I(N__45421));
    InMux I__9707 (
            .O(N__45424),
            .I(N__45418));
    Span4Mux_h I__9706 (
            .O(N__45421),
            .I(N__45415));
    LocalMux I__9705 (
            .O(N__45418),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__9704 (
            .O(N__45415),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__9703 (
            .O(N__45410),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__9702 (
            .O(N__45407),
            .I(N__45369));
    InMux I__9701 (
            .O(N__45406),
            .I(N__45369));
    InMux I__9700 (
            .O(N__45405),
            .I(N__45369));
    InMux I__9699 (
            .O(N__45404),
            .I(N__45369));
    InMux I__9698 (
            .O(N__45403),
            .I(N__45364));
    InMux I__9697 (
            .O(N__45402),
            .I(N__45364));
    InMux I__9696 (
            .O(N__45401),
            .I(N__45355));
    InMux I__9695 (
            .O(N__45400),
            .I(N__45355));
    InMux I__9694 (
            .O(N__45399),
            .I(N__45355));
    InMux I__9693 (
            .O(N__45398),
            .I(N__45355));
    InMux I__9692 (
            .O(N__45397),
            .I(N__45346));
    InMux I__9691 (
            .O(N__45396),
            .I(N__45346));
    InMux I__9690 (
            .O(N__45395),
            .I(N__45346));
    InMux I__9689 (
            .O(N__45394),
            .I(N__45346));
    InMux I__9688 (
            .O(N__45393),
            .I(N__45337));
    InMux I__9687 (
            .O(N__45392),
            .I(N__45337));
    InMux I__9686 (
            .O(N__45391),
            .I(N__45337));
    InMux I__9685 (
            .O(N__45390),
            .I(N__45337));
    InMux I__9684 (
            .O(N__45389),
            .I(N__45328));
    InMux I__9683 (
            .O(N__45388),
            .I(N__45328));
    InMux I__9682 (
            .O(N__45387),
            .I(N__45328));
    InMux I__9681 (
            .O(N__45386),
            .I(N__45328));
    InMux I__9680 (
            .O(N__45385),
            .I(N__45319));
    InMux I__9679 (
            .O(N__45384),
            .I(N__45319));
    InMux I__9678 (
            .O(N__45383),
            .I(N__45319));
    InMux I__9677 (
            .O(N__45382),
            .I(N__45319));
    InMux I__9676 (
            .O(N__45381),
            .I(N__45310));
    InMux I__9675 (
            .O(N__45380),
            .I(N__45310));
    InMux I__9674 (
            .O(N__45379),
            .I(N__45310));
    InMux I__9673 (
            .O(N__45378),
            .I(N__45310));
    LocalMux I__9672 (
            .O(N__45369),
            .I(N__45303));
    LocalMux I__9671 (
            .O(N__45364),
            .I(N__45303));
    LocalMux I__9670 (
            .O(N__45355),
            .I(N__45303));
    LocalMux I__9669 (
            .O(N__45346),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__9668 (
            .O(N__45337),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__9667 (
            .O(N__45328),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__9666 (
            .O(N__45319),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__9665 (
            .O(N__45310),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__9664 (
            .O(N__45303),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__9663 (
            .O(N__45290),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CascadeMux I__9662 (
            .O(N__45287),
            .I(N__45284));
    InMux I__9661 (
            .O(N__45284),
            .I(N__45280));
    InMux I__9660 (
            .O(N__45283),
            .I(N__45277));
    LocalMux I__9659 (
            .O(N__45280),
            .I(N__45274));
    LocalMux I__9658 (
            .O(N__45277),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv12 I__9657 (
            .O(N__45274),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CEMux I__9656 (
            .O(N__45269),
            .I(N__45264));
    CEMux I__9655 (
            .O(N__45268),
            .I(N__45261));
    CEMux I__9654 (
            .O(N__45267),
            .I(N__45258));
    LocalMux I__9653 (
            .O(N__45264),
            .I(N__45255));
    LocalMux I__9652 (
            .O(N__45261),
            .I(N__45252));
    LocalMux I__9651 (
            .O(N__45258),
            .I(N__45248));
    Span4Mux_v I__9650 (
            .O(N__45255),
            .I(N__45243));
    Span4Mux_v I__9649 (
            .O(N__45252),
            .I(N__45243));
    CEMux I__9648 (
            .O(N__45251),
            .I(N__45240));
    Span4Mux_v I__9647 (
            .O(N__45248),
            .I(N__45233));
    Span4Mux_h I__9646 (
            .O(N__45243),
            .I(N__45233));
    LocalMux I__9645 (
            .O(N__45240),
            .I(N__45233));
    Span4Mux_h I__9644 (
            .O(N__45233),
            .I(N__45230));
    Odrv4 I__9643 (
            .O(N__45230),
            .I(\delay_measurement_inst.delay_hc_timer.N_166_i ));
    InMux I__9642 (
            .O(N__45227),
            .I(N__45224));
    LocalMux I__9641 (
            .O(N__45224),
            .I(N__45220));
    CascadeMux I__9640 (
            .O(N__45223),
            .I(N__45217));
    Span4Mux_h I__9639 (
            .O(N__45220),
            .I(N__45213));
    InMux I__9638 (
            .O(N__45217),
            .I(N__45210));
    InMux I__9637 (
            .O(N__45216),
            .I(N__45207));
    Span4Mux_v I__9636 (
            .O(N__45213),
            .I(N__45202));
    LocalMux I__9635 (
            .O(N__45210),
            .I(N__45202));
    LocalMux I__9634 (
            .O(N__45207),
            .I(N__45197));
    Span4Mux_v I__9633 (
            .O(N__45202),
            .I(N__45197));
    Odrv4 I__9632 (
            .O(N__45197),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__9631 (
            .O(N__45194),
            .I(bfn_17_11_0_));
    InMux I__9630 (
            .O(N__45191),
            .I(N__45187));
    CascadeMux I__9629 (
            .O(N__45190),
            .I(N__45184));
    LocalMux I__9628 (
            .O(N__45187),
            .I(N__45181));
    InMux I__9627 (
            .O(N__45184),
            .I(N__45177));
    Span4Mux_h I__9626 (
            .O(N__45181),
            .I(N__45174));
    InMux I__9625 (
            .O(N__45180),
            .I(N__45171));
    LocalMux I__9624 (
            .O(N__45177),
            .I(N__45168));
    Span4Mux_v I__9623 (
            .O(N__45174),
            .I(N__45165));
    LocalMux I__9622 (
            .O(N__45171),
            .I(N__45160));
    Span4Mux_v I__9621 (
            .O(N__45168),
            .I(N__45160));
    Odrv4 I__9620 (
            .O(N__45165),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__9619 (
            .O(N__45160),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__9618 (
            .O(N__45155),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__9617 (
            .O(N__45152),
            .I(N__45146));
    InMux I__9616 (
            .O(N__45151),
            .I(N__45146));
    LocalMux I__9615 (
            .O(N__45146),
            .I(N__45142));
    InMux I__9614 (
            .O(N__45145),
            .I(N__45139));
    Span4Mux_h I__9613 (
            .O(N__45142),
            .I(N__45136));
    LocalMux I__9612 (
            .O(N__45139),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv4 I__9611 (
            .O(N__45136),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__9610 (
            .O(N__45131),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__9609 (
            .O(N__45128),
            .I(N__45122));
    InMux I__9608 (
            .O(N__45127),
            .I(N__45122));
    LocalMux I__9607 (
            .O(N__45122),
            .I(N__45118));
    InMux I__9606 (
            .O(N__45121),
            .I(N__45115));
    Span4Mux_h I__9605 (
            .O(N__45118),
            .I(N__45112));
    LocalMux I__9604 (
            .O(N__45115),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__9603 (
            .O(N__45112),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__9602 (
            .O(N__45107),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__9601 (
            .O(N__45104),
            .I(N__45100));
    CascadeMux I__9600 (
            .O(N__45103),
            .I(N__45097));
    InMux I__9599 (
            .O(N__45100),
            .I(N__45092));
    InMux I__9598 (
            .O(N__45097),
            .I(N__45092));
    LocalMux I__9597 (
            .O(N__45092),
            .I(N__45088));
    InMux I__9596 (
            .O(N__45091),
            .I(N__45085));
    Span4Mux_h I__9595 (
            .O(N__45088),
            .I(N__45082));
    LocalMux I__9594 (
            .O(N__45085),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__9593 (
            .O(N__45082),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__9592 (
            .O(N__45077),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__9591 (
            .O(N__45074),
            .I(N__45070));
    CascadeMux I__9590 (
            .O(N__45073),
            .I(N__45067));
    InMux I__9589 (
            .O(N__45070),
            .I(N__45062));
    InMux I__9588 (
            .O(N__45067),
            .I(N__45062));
    LocalMux I__9587 (
            .O(N__45062),
            .I(N__45058));
    InMux I__9586 (
            .O(N__45061),
            .I(N__45055));
    Span4Mux_h I__9585 (
            .O(N__45058),
            .I(N__45052));
    LocalMux I__9584 (
            .O(N__45055),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__9583 (
            .O(N__45052),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__9582 (
            .O(N__45047),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__9581 (
            .O(N__45044),
            .I(N__45041));
    InMux I__9580 (
            .O(N__45041),
            .I(N__45037));
    InMux I__9579 (
            .O(N__45040),
            .I(N__45034));
    LocalMux I__9578 (
            .O(N__45037),
            .I(N__45028));
    LocalMux I__9577 (
            .O(N__45034),
            .I(N__45028));
    InMux I__9576 (
            .O(N__45033),
            .I(N__45025));
    Span4Mux_h I__9575 (
            .O(N__45028),
            .I(N__45022));
    LocalMux I__9574 (
            .O(N__45025),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__9573 (
            .O(N__45022),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__9572 (
            .O(N__45017),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    CascadeMux I__9571 (
            .O(N__45014),
            .I(N__45010));
    CascadeMux I__9570 (
            .O(N__45013),
            .I(N__45007));
    InMux I__9569 (
            .O(N__45010),
            .I(N__45001));
    InMux I__9568 (
            .O(N__45007),
            .I(N__45001));
    InMux I__9567 (
            .O(N__45006),
            .I(N__44998));
    LocalMux I__9566 (
            .O(N__45001),
            .I(N__44995));
    LocalMux I__9565 (
            .O(N__44998),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv12 I__9564 (
            .O(N__44995),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__9563 (
            .O(N__44990),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__9562 (
            .O(N__44987),
            .I(N__44983));
    CascadeMux I__9561 (
            .O(N__44986),
            .I(N__44980));
    InMux I__9560 (
            .O(N__44983),
            .I(N__44974));
    InMux I__9559 (
            .O(N__44980),
            .I(N__44974));
    InMux I__9558 (
            .O(N__44979),
            .I(N__44971));
    LocalMux I__9557 (
            .O(N__44974),
            .I(N__44968));
    LocalMux I__9556 (
            .O(N__44971),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv12 I__9555 (
            .O(N__44968),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__9554 (
            .O(N__44963),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    CascadeMux I__9553 (
            .O(N__44960),
            .I(N__44957));
    InMux I__9552 (
            .O(N__44957),
            .I(N__44952));
    InMux I__9551 (
            .O(N__44956),
            .I(N__44949));
    InMux I__9550 (
            .O(N__44955),
            .I(N__44946));
    LocalMux I__9549 (
            .O(N__44952),
            .I(N__44941));
    LocalMux I__9548 (
            .O(N__44949),
            .I(N__44941));
    LocalMux I__9547 (
            .O(N__44946),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv12 I__9546 (
            .O(N__44941),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__9545 (
            .O(N__44936),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    CascadeMux I__9544 (
            .O(N__44933),
            .I(N__44930));
    InMux I__9543 (
            .O(N__44930),
            .I(N__44925));
    InMux I__9542 (
            .O(N__44929),
            .I(N__44922));
    InMux I__9541 (
            .O(N__44928),
            .I(N__44919));
    LocalMux I__9540 (
            .O(N__44925),
            .I(N__44914));
    LocalMux I__9539 (
            .O(N__44922),
            .I(N__44914));
    LocalMux I__9538 (
            .O(N__44919),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv12 I__9537 (
            .O(N__44914),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__9536 (
            .O(N__44909),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__9535 (
            .O(N__44906),
            .I(N__44903));
    InMux I__9534 (
            .O(N__44903),
            .I(N__44900));
    LocalMux I__9533 (
            .O(N__44900),
            .I(N__44895));
    InMux I__9532 (
            .O(N__44899),
            .I(N__44892));
    InMux I__9531 (
            .O(N__44898),
            .I(N__44889));
    Span4Mux_h I__9530 (
            .O(N__44895),
            .I(N__44886));
    LocalMux I__9529 (
            .O(N__44892),
            .I(N__44883));
    LocalMux I__9528 (
            .O(N__44889),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__9527 (
            .O(N__44886),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv12 I__9526 (
            .O(N__44883),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__9525 (
            .O(N__44876),
            .I(bfn_17_10_0_));
    CascadeMux I__9524 (
            .O(N__44873),
            .I(N__44870));
    InMux I__9523 (
            .O(N__44870),
            .I(N__44867));
    LocalMux I__9522 (
            .O(N__44867),
            .I(N__44862));
    InMux I__9521 (
            .O(N__44866),
            .I(N__44859));
    InMux I__9520 (
            .O(N__44865),
            .I(N__44856));
    Span4Mux_h I__9519 (
            .O(N__44862),
            .I(N__44853));
    LocalMux I__9518 (
            .O(N__44859),
            .I(N__44850));
    LocalMux I__9517 (
            .O(N__44856),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__9516 (
            .O(N__44853),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv12 I__9515 (
            .O(N__44850),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__9514 (
            .O(N__44843),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__9513 (
            .O(N__44840),
            .I(N__44833));
    InMux I__9512 (
            .O(N__44839),
            .I(N__44833));
    InMux I__9511 (
            .O(N__44838),
            .I(N__44830));
    LocalMux I__9510 (
            .O(N__44833),
            .I(N__44827));
    LocalMux I__9509 (
            .O(N__44830),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv12 I__9508 (
            .O(N__44827),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__9507 (
            .O(N__44822),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__9506 (
            .O(N__44819),
            .I(N__44812));
    InMux I__9505 (
            .O(N__44818),
            .I(N__44812));
    InMux I__9504 (
            .O(N__44817),
            .I(N__44809));
    LocalMux I__9503 (
            .O(N__44812),
            .I(N__44806));
    LocalMux I__9502 (
            .O(N__44809),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv12 I__9501 (
            .O(N__44806),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__9500 (
            .O(N__44801),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    CascadeMux I__9499 (
            .O(N__44798),
            .I(N__44795));
    InMux I__9498 (
            .O(N__44795),
            .I(N__44791));
    InMux I__9497 (
            .O(N__44794),
            .I(N__44788));
    LocalMux I__9496 (
            .O(N__44791),
            .I(N__44785));
    LocalMux I__9495 (
            .O(N__44788),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv12 I__9494 (
            .O(N__44785),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__9493 (
            .O(N__44780),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    CascadeMux I__9492 (
            .O(N__44777),
            .I(N__44773));
    CascadeMux I__9491 (
            .O(N__44776),
            .I(N__44770));
    InMux I__9490 (
            .O(N__44773),
            .I(N__44765));
    InMux I__9489 (
            .O(N__44770),
            .I(N__44765));
    LocalMux I__9488 (
            .O(N__44765),
            .I(N__44761));
    InMux I__9487 (
            .O(N__44764),
            .I(N__44758));
    Span4Mux_h I__9486 (
            .O(N__44761),
            .I(N__44755));
    LocalMux I__9485 (
            .O(N__44758),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__9484 (
            .O(N__44755),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__9483 (
            .O(N__44750),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__9482 (
            .O(N__44747),
            .I(N__44743));
    CascadeMux I__9481 (
            .O(N__44746),
            .I(N__44740));
    InMux I__9480 (
            .O(N__44743),
            .I(N__44735));
    InMux I__9479 (
            .O(N__44740),
            .I(N__44735));
    LocalMux I__9478 (
            .O(N__44735),
            .I(N__44731));
    InMux I__9477 (
            .O(N__44734),
            .I(N__44728));
    Span4Mux_h I__9476 (
            .O(N__44731),
            .I(N__44725));
    LocalMux I__9475 (
            .O(N__44728),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__9474 (
            .O(N__44725),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__9473 (
            .O(N__44720),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    CascadeMux I__9472 (
            .O(N__44717),
            .I(N__44714));
    InMux I__9471 (
            .O(N__44714),
            .I(N__44710));
    InMux I__9470 (
            .O(N__44713),
            .I(N__44707));
    LocalMux I__9469 (
            .O(N__44710),
            .I(N__44701));
    LocalMux I__9468 (
            .O(N__44707),
            .I(N__44701));
    InMux I__9467 (
            .O(N__44706),
            .I(N__44698));
    Span4Mux_v I__9466 (
            .O(N__44701),
            .I(N__44695));
    LocalMux I__9465 (
            .O(N__44698),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__9464 (
            .O(N__44695),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__9463 (
            .O(N__44690),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__9462 (
            .O(N__44687),
            .I(N__44681));
    InMux I__9461 (
            .O(N__44686),
            .I(N__44681));
    LocalMux I__9460 (
            .O(N__44681),
            .I(N__44677));
    InMux I__9459 (
            .O(N__44680),
            .I(N__44674));
    Span4Mux_v I__9458 (
            .O(N__44677),
            .I(N__44671));
    LocalMux I__9457 (
            .O(N__44674),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__9456 (
            .O(N__44671),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__9455 (
            .O(N__44666),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__9454 (
            .O(N__44663),
            .I(N__44660));
    InMux I__9453 (
            .O(N__44660),
            .I(N__44657));
    LocalMux I__9452 (
            .O(N__44657),
            .I(N__44652));
    InMux I__9451 (
            .O(N__44656),
            .I(N__44649));
    InMux I__9450 (
            .O(N__44655),
            .I(N__44646));
    Span4Mux_h I__9449 (
            .O(N__44652),
            .I(N__44643));
    LocalMux I__9448 (
            .O(N__44649),
            .I(N__44640));
    LocalMux I__9447 (
            .O(N__44646),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__9446 (
            .O(N__44643),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv12 I__9445 (
            .O(N__44640),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__9444 (
            .O(N__44633),
            .I(bfn_17_9_0_));
    CascadeMux I__9443 (
            .O(N__44630),
            .I(N__44627));
    InMux I__9442 (
            .O(N__44627),
            .I(N__44623));
    CascadeMux I__9441 (
            .O(N__44626),
            .I(N__44620));
    LocalMux I__9440 (
            .O(N__44623),
            .I(N__44616));
    InMux I__9439 (
            .O(N__44620),
            .I(N__44613));
    InMux I__9438 (
            .O(N__44619),
            .I(N__44610));
    Span4Mux_h I__9437 (
            .O(N__44616),
            .I(N__44607));
    LocalMux I__9436 (
            .O(N__44613),
            .I(N__44604));
    LocalMux I__9435 (
            .O(N__44610),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__9434 (
            .O(N__44607),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv12 I__9433 (
            .O(N__44604),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__9432 (
            .O(N__44597),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__9431 (
            .O(N__44594),
            .I(N__44588));
    InMux I__9430 (
            .O(N__44593),
            .I(N__44588));
    LocalMux I__9429 (
            .O(N__44588),
            .I(N__44584));
    InMux I__9428 (
            .O(N__44587),
            .I(N__44581));
    Span4Mux_h I__9427 (
            .O(N__44584),
            .I(N__44578));
    LocalMux I__9426 (
            .O(N__44581),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__9425 (
            .O(N__44578),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__9424 (
            .O(N__44573),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__9423 (
            .O(N__44570),
            .I(N__44564));
    InMux I__9422 (
            .O(N__44569),
            .I(N__44564));
    LocalMux I__9421 (
            .O(N__44564),
            .I(N__44560));
    InMux I__9420 (
            .O(N__44563),
            .I(N__44557));
    Span4Mux_h I__9419 (
            .O(N__44560),
            .I(N__44554));
    LocalMux I__9418 (
            .O(N__44557),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv4 I__9417 (
            .O(N__44554),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__9416 (
            .O(N__44549),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__9415 (
            .O(N__44546),
            .I(N__44540));
    InMux I__9414 (
            .O(N__44545),
            .I(N__44540));
    LocalMux I__9413 (
            .O(N__44540),
            .I(N__44536));
    InMux I__9412 (
            .O(N__44539),
            .I(N__44533));
    Span4Mux_s2_v I__9411 (
            .O(N__44536),
            .I(N__44530));
    LocalMux I__9410 (
            .O(N__44533),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__9409 (
            .O(N__44530),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__9408 (
            .O(N__44525),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__9407 (
            .O(N__44522),
            .I(N__44518));
    CascadeMux I__9406 (
            .O(N__44521),
            .I(N__44515));
    InMux I__9405 (
            .O(N__44518),
            .I(N__44510));
    InMux I__9404 (
            .O(N__44515),
            .I(N__44510));
    LocalMux I__9403 (
            .O(N__44510),
            .I(N__44506));
    InMux I__9402 (
            .O(N__44509),
            .I(N__44503));
    Span4Mux_s2_v I__9401 (
            .O(N__44506),
            .I(N__44500));
    LocalMux I__9400 (
            .O(N__44503),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__9399 (
            .O(N__44500),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__9398 (
            .O(N__44495),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__9397 (
            .O(N__44492),
            .I(N__44488));
    CascadeMux I__9396 (
            .O(N__44491),
            .I(N__44485));
    InMux I__9395 (
            .O(N__44488),
            .I(N__44480));
    InMux I__9394 (
            .O(N__44485),
            .I(N__44480));
    LocalMux I__9393 (
            .O(N__44480),
            .I(N__44476));
    InMux I__9392 (
            .O(N__44479),
            .I(N__44473));
    Span4Mux_s2_v I__9391 (
            .O(N__44476),
            .I(N__44470));
    LocalMux I__9390 (
            .O(N__44473),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__9389 (
            .O(N__44470),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__9388 (
            .O(N__44465),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    CascadeMux I__9387 (
            .O(N__44462),
            .I(N__44459));
    InMux I__9386 (
            .O(N__44459),
            .I(N__44455));
    InMux I__9385 (
            .O(N__44458),
            .I(N__44452));
    LocalMux I__9384 (
            .O(N__44455),
            .I(N__44446));
    LocalMux I__9383 (
            .O(N__44452),
            .I(N__44446));
    InMux I__9382 (
            .O(N__44451),
            .I(N__44443));
    Span4Mux_s3_v I__9381 (
            .O(N__44446),
            .I(N__44440));
    LocalMux I__9380 (
            .O(N__44443),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__9379 (
            .O(N__44440),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__9378 (
            .O(N__44435),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    CascadeMux I__9377 (
            .O(N__44432),
            .I(N__44429));
    InMux I__9376 (
            .O(N__44429),
            .I(N__44425));
    InMux I__9375 (
            .O(N__44428),
            .I(N__44422));
    LocalMux I__9374 (
            .O(N__44425),
            .I(N__44416));
    LocalMux I__9373 (
            .O(N__44422),
            .I(N__44416));
    InMux I__9372 (
            .O(N__44421),
            .I(N__44413));
    Span4Mux_s3_v I__9371 (
            .O(N__44416),
            .I(N__44410));
    LocalMux I__9370 (
            .O(N__44413),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__9369 (
            .O(N__44410),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__9368 (
            .O(N__44405),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__9367 (
            .O(N__44402),
            .I(N__44399));
    InMux I__9366 (
            .O(N__44399),
            .I(N__44396));
    LocalMux I__9365 (
            .O(N__44396),
            .I(N__44391));
    InMux I__9364 (
            .O(N__44395),
            .I(N__44388));
    InMux I__9363 (
            .O(N__44394),
            .I(N__44385));
    Span4Mux_h I__9362 (
            .O(N__44391),
            .I(N__44382));
    LocalMux I__9361 (
            .O(N__44388),
            .I(N__44379));
    LocalMux I__9360 (
            .O(N__44385),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__9359 (
            .O(N__44382),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv12 I__9358 (
            .O(N__44379),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__9357 (
            .O(N__44372),
            .I(bfn_17_8_0_));
    CascadeMux I__9356 (
            .O(N__44369),
            .I(N__44366));
    InMux I__9355 (
            .O(N__44366),
            .I(N__44363));
    LocalMux I__9354 (
            .O(N__44363),
            .I(N__44358));
    InMux I__9353 (
            .O(N__44362),
            .I(N__44355));
    InMux I__9352 (
            .O(N__44361),
            .I(N__44352));
    Sp12to4 I__9351 (
            .O(N__44358),
            .I(N__44347));
    LocalMux I__9350 (
            .O(N__44355),
            .I(N__44347));
    LocalMux I__9349 (
            .O(N__44352),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv12 I__9348 (
            .O(N__44347),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__9347 (
            .O(N__44342),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__9346 (
            .O(N__44339),
            .I(N__44333));
    InMux I__9345 (
            .O(N__44338),
            .I(N__44333));
    LocalMux I__9344 (
            .O(N__44333),
            .I(N__44329));
    InMux I__9343 (
            .O(N__44332),
            .I(N__44326));
    Span4Mux_h I__9342 (
            .O(N__44329),
            .I(N__44323));
    LocalMux I__9341 (
            .O(N__44326),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__9340 (
            .O(N__44323),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__9339 (
            .O(N__44318),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__9338 (
            .O(N__44315),
            .I(N__44309));
    InMux I__9337 (
            .O(N__44314),
            .I(N__44309));
    LocalMux I__9336 (
            .O(N__44309),
            .I(N__44305));
    InMux I__9335 (
            .O(N__44308),
            .I(N__44302));
    Span4Mux_h I__9334 (
            .O(N__44305),
            .I(N__44299));
    LocalMux I__9333 (
            .O(N__44302),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__9332 (
            .O(N__44299),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__9331 (
            .O(N__44294),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__9330 (
            .O(N__44291),
            .I(N__44288));
    LocalMux I__9329 (
            .O(N__44288),
            .I(N__44285));
    Span4Mux_h I__9328 (
            .O(N__44285),
            .I(N__44281));
    InMux I__9327 (
            .O(N__44284),
            .I(N__44278));
    Odrv4 I__9326 (
            .O(N__44281),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    LocalMux I__9325 (
            .O(N__44278),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__9324 (
            .O(N__44273),
            .I(bfn_17_6_0_));
    InMux I__9323 (
            .O(N__44270),
            .I(N__44267));
    LocalMux I__9322 (
            .O(N__44267),
            .I(N__44264));
    Span4Mux_v I__9321 (
            .O(N__44264),
            .I(N__44260));
    InMux I__9320 (
            .O(N__44263),
            .I(N__44257));
    Odrv4 I__9319 (
            .O(N__44260),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    LocalMux I__9318 (
            .O(N__44257),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__9317 (
            .O(N__44252),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__9316 (
            .O(N__44249),
            .I(N__44245));
    InMux I__9315 (
            .O(N__44248),
            .I(N__44242));
    LocalMux I__9314 (
            .O(N__44245),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__9313 (
            .O(N__44242),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__9312 (
            .O(N__44237),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__9311 (
            .O(N__44234),
            .I(N__44231));
    LocalMux I__9310 (
            .O(N__44231),
            .I(N__44227));
    InMux I__9309 (
            .O(N__44230),
            .I(N__44224));
    Odrv4 I__9308 (
            .O(N__44227),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__9307 (
            .O(N__44224),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__9306 (
            .O(N__44219),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__9305 (
            .O(N__44216),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__9304 (
            .O(N__44213),
            .I(N__44210));
    LocalMux I__9303 (
            .O(N__44210),
            .I(N__44206));
    InMux I__9302 (
            .O(N__44209),
            .I(N__44203));
    Span4Mux_h I__9301 (
            .O(N__44206),
            .I(N__44198));
    LocalMux I__9300 (
            .O(N__44203),
            .I(N__44198));
    Odrv4 I__9299 (
            .O(N__44198),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    CEMux I__9298 (
            .O(N__44195),
            .I(N__44189));
    CEMux I__9297 (
            .O(N__44194),
            .I(N__44186));
    CEMux I__9296 (
            .O(N__44193),
            .I(N__44183));
    CEMux I__9295 (
            .O(N__44192),
            .I(N__44179));
    LocalMux I__9294 (
            .O(N__44189),
            .I(N__44176));
    LocalMux I__9293 (
            .O(N__44186),
            .I(N__44171));
    LocalMux I__9292 (
            .O(N__44183),
            .I(N__44171));
    CEMux I__9291 (
            .O(N__44182),
            .I(N__44168));
    LocalMux I__9290 (
            .O(N__44179),
            .I(N__44165));
    Span4Mux_v I__9289 (
            .O(N__44176),
            .I(N__44158));
    Span4Mux_v I__9288 (
            .O(N__44171),
            .I(N__44158));
    LocalMux I__9287 (
            .O(N__44168),
            .I(N__44158));
    Span4Mux_v I__9286 (
            .O(N__44165),
            .I(N__44153));
    Span4Mux_h I__9285 (
            .O(N__44158),
            .I(N__44153));
    Odrv4 I__9284 (
            .O(N__44153),
            .I(\delay_measurement_inst.delay_hc_timer.N_165_i ));
    InMux I__9283 (
            .O(N__44150),
            .I(N__44146));
    InMux I__9282 (
            .O(N__44149),
            .I(N__44143));
    LocalMux I__9281 (
            .O(N__44146),
            .I(N__44139));
    LocalMux I__9280 (
            .O(N__44143),
            .I(N__44136));
    InMux I__9279 (
            .O(N__44142),
            .I(N__44133));
    Odrv4 I__9278 (
            .O(N__44139),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv12 I__9277 (
            .O(N__44136),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__9276 (
            .O(N__44133),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__9275 (
            .O(N__44126),
            .I(bfn_17_7_0_));
    CascadeMux I__9274 (
            .O(N__44123),
            .I(N__44120));
    InMux I__9273 (
            .O(N__44120),
            .I(N__44116));
    InMux I__9272 (
            .O(N__44119),
            .I(N__44112));
    LocalMux I__9271 (
            .O(N__44116),
            .I(N__44109));
    InMux I__9270 (
            .O(N__44115),
            .I(N__44106));
    LocalMux I__9269 (
            .O(N__44112),
            .I(N__44101));
    Span4Mux_s2_v I__9268 (
            .O(N__44109),
            .I(N__44101));
    LocalMux I__9267 (
            .O(N__44106),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__9266 (
            .O(N__44101),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__9265 (
            .O(N__44096),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    CascadeMux I__9264 (
            .O(N__44093),
            .I(N__44089));
    InMux I__9263 (
            .O(N__44092),
            .I(N__44086));
    InMux I__9262 (
            .O(N__44089),
            .I(N__44083));
    LocalMux I__9261 (
            .O(N__44086),
            .I(N__44077));
    LocalMux I__9260 (
            .O(N__44083),
            .I(N__44077));
    InMux I__9259 (
            .O(N__44082),
            .I(N__44074));
    Span4Mux_s2_v I__9258 (
            .O(N__44077),
            .I(N__44071));
    LocalMux I__9257 (
            .O(N__44074),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__9256 (
            .O(N__44071),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__9255 (
            .O(N__44066),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__9254 (
            .O(N__44063),
            .I(N__44060));
    LocalMux I__9253 (
            .O(N__44060),
            .I(N__44057));
    Span4Mux_h I__9252 (
            .O(N__44057),
            .I(N__44053));
    InMux I__9251 (
            .O(N__44056),
            .I(N__44050));
    Odrv4 I__9250 (
            .O(N__44053),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    LocalMux I__9249 (
            .O(N__44050),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__9248 (
            .O(N__44045),
            .I(bfn_17_5_0_));
    InMux I__9247 (
            .O(N__44042),
            .I(N__44039));
    LocalMux I__9246 (
            .O(N__44039),
            .I(N__44036));
    Span4Mux_h I__9245 (
            .O(N__44036),
            .I(N__44032));
    InMux I__9244 (
            .O(N__44035),
            .I(N__44029));
    Odrv4 I__9243 (
            .O(N__44032),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__9242 (
            .O(N__44029),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__9241 (
            .O(N__44024),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__9240 (
            .O(N__44021),
            .I(N__44018));
    LocalMux I__9239 (
            .O(N__44018),
            .I(N__44015));
    Span4Mux_v I__9238 (
            .O(N__44015),
            .I(N__44011));
    InMux I__9237 (
            .O(N__44014),
            .I(N__44008));
    Odrv4 I__9236 (
            .O(N__44011),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__9235 (
            .O(N__44008),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__9234 (
            .O(N__44003),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__9233 (
            .O(N__44000),
            .I(N__43996));
    CascadeMux I__9232 (
            .O(N__43999),
            .I(N__43993));
    LocalMux I__9231 (
            .O(N__43996),
            .I(N__43990));
    InMux I__9230 (
            .O(N__43993),
            .I(N__43987));
    Odrv4 I__9229 (
            .O(N__43990),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__9228 (
            .O(N__43987),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__9227 (
            .O(N__43982),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__9226 (
            .O(N__43979),
            .I(N__43976));
    LocalMux I__9225 (
            .O(N__43976),
            .I(N__43972));
    CascadeMux I__9224 (
            .O(N__43975),
            .I(N__43969));
    Span4Mux_h I__9223 (
            .O(N__43972),
            .I(N__43966));
    InMux I__9222 (
            .O(N__43969),
            .I(N__43963));
    Odrv4 I__9221 (
            .O(N__43966),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__9220 (
            .O(N__43963),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__9219 (
            .O(N__43958),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__9218 (
            .O(N__43955),
            .I(N__43952));
    LocalMux I__9217 (
            .O(N__43952),
            .I(N__43949));
    Span4Mux_h I__9216 (
            .O(N__43949),
            .I(N__43945));
    InMux I__9215 (
            .O(N__43948),
            .I(N__43942));
    Odrv4 I__9214 (
            .O(N__43945),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__9213 (
            .O(N__43942),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__9212 (
            .O(N__43937),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__9211 (
            .O(N__43934),
            .I(N__43931));
    LocalMux I__9210 (
            .O(N__43931),
            .I(N__43927));
    CascadeMux I__9209 (
            .O(N__43930),
            .I(N__43924));
    Span4Mux_v I__9208 (
            .O(N__43927),
            .I(N__43921));
    InMux I__9207 (
            .O(N__43924),
            .I(N__43918));
    Odrv4 I__9206 (
            .O(N__43921),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__9205 (
            .O(N__43918),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__9204 (
            .O(N__43913),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__9203 (
            .O(N__43910),
            .I(N__43907));
    LocalMux I__9202 (
            .O(N__43907),
            .I(N__43904));
    Span4Mux_h I__9201 (
            .O(N__43904),
            .I(N__43900));
    InMux I__9200 (
            .O(N__43903),
            .I(N__43897));
    Odrv4 I__9199 (
            .O(N__43900),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__9198 (
            .O(N__43897),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__9197 (
            .O(N__43892),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__9196 (
            .O(N__43889),
            .I(N__43886));
    LocalMux I__9195 (
            .O(N__43886),
            .I(N__43882));
    InMux I__9194 (
            .O(N__43885),
            .I(N__43879));
    Span4Mux_h I__9193 (
            .O(N__43882),
            .I(N__43876));
    LocalMux I__9192 (
            .O(N__43879),
            .I(N__43873));
    Odrv4 I__9191 (
            .O(N__43876),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    Odrv4 I__9190 (
            .O(N__43873),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__9189 (
            .O(N__43868),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__9188 (
            .O(N__43865),
            .I(N__43862));
    LocalMux I__9187 (
            .O(N__43862),
            .I(N__43859));
    Span4Mux_h I__9186 (
            .O(N__43859),
            .I(N__43855));
    InMux I__9185 (
            .O(N__43858),
            .I(N__43852));
    Odrv4 I__9184 (
            .O(N__43855),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__9183 (
            .O(N__43852),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__9182 (
            .O(N__43847),
            .I(bfn_17_4_0_));
    InMux I__9181 (
            .O(N__43844),
            .I(N__43841));
    LocalMux I__9180 (
            .O(N__43841),
            .I(N__43838));
    Span4Mux_v I__9179 (
            .O(N__43838),
            .I(N__43834));
    InMux I__9178 (
            .O(N__43837),
            .I(N__43831));
    Odrv4 I__9177 (
            .O(N__43834),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__9176 (
            .O(N__43831),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__9175 (
            .O(N__43826),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__9174 (
            .O(N__43823),
            .I(N__43820));
    LocalMux I__9173 (
            .O(N__43820),
            .I(N__43817));
    Span4Mux_h I__9172 (
            .O(N__43817),
            .I(N__43813));
    InMux I__9171 (
            .O(N__43816),
            .I(N__43810));
    Odrv4 I__9170 (
            .O(N__43813),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__9169 (
            .O(N__43810),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__9168 (
            .O(N__43805),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__9167 (
            .O(N__43802),
            .I(N__43799));
    LocalMux I__9166 (
            .O(N__43799),
            .I(N__43796));
    Span4Mux_h I__9165 (
            .O(N__43796),
            .I(N__43792));
    InMux I__9164 (
            .O(N__43795),
            .I(N__43789));
    Odrv4 I__9163 (
            .O(N__43792),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    LocalMux I__9162 (
            .O(N__43789),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__9161 (
            .O(N__43784),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__9160 (
            .O(N__43781),
            .I(N__43778));
    LocalMux I__9159 (
            .O(N__43778),
            .I(N__43775));
    Span4Mux_h I__9158 (
            .O(N__43775),
            .I(N__43771));
    InMux I__9157 (
            .O(N__43774),
            .I(N__43768));
    Odrv4 I__9156 (
            .O(N__43771),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    LocalMux I__9155 (
            .O(N__43768),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__9154 (
            .O(N__43763),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__9153 (
            .O(N__43760),
            .I(N__43757));
    LocalMux I__9152 (
            .O(N__43757),
            .I(N__43753));
    InMux I__9151 (
            .O(N__43756),
            .I(N__43750));
    Odrv4 I__9150 (
            .O(N__43753),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__9149 (
            .O(N__43750),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__9148 (
            .O(N__43745),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__9147 (
            .O(N__43742),
            .I(N__43739));
    LocalMux I__9146 (
            .O(N__43739),
            .I(N__43736));
    Span4Mux_v I__9145 (
            .O(N__43736),
            .I(N__43733));
    Span4Mux_h I__9144 (
            .O(N__43733),
            .I(N__43729));
    InMux I__9143 (
            .O(N__43732),
            .I(N__43726));
    Odrv4 I__9142 (
            .O(N__43729),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__9141 (
            .O(N__43726),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__9140 (
            .O(N__43721),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__9139 (
            .O(N__43718),
            .I(N__43715));
    LocalMux I__9138 (
            .O(N__43715),
            .I(N__43711));
    CascadeMux I__9137 (
            .O(N__43714),
            .I(N__43708));
    Span4Mux_v I__9136 (
            .O(N__43711),
            .I(N__43705));
    InMux I__9135 (
            .O(N__43708),
            .I(N__43702));
    Odrv4 I__9134 (
            .O(N__43705),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__9133 (
            .O(N__43702),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__9132 (
            .O(N__43697),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__9131 (
            .O(N__43694),
            .I(N__43691));
    LocalMux I__9130 (
            .O(N__43691),
            .I(N__43688));
    Span4Mux_v I__9129 (
            .O(N__43688),
            .I(N__43684));
    InMux I__9128 (
            .O(N__43687),
            .I(N__43681));
    Odrv4 I__9127 (
            .O(N__43684),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__9126 (
            .O(N__43681),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__9125 (
            .O(N__43676),
            .I(N__43673));
    LocalMux I__9124 (
            .O(N__43673),
            .I(N__43670));
    Span4Mux_v I__9123 (
            .O(N__43670),
            .I(N__43666));
    InMux I__9122 (
            .O(N__43669),
            .I(N__43663));
    Odrv4 I__9121 (
            .O(N__43666),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__9120 (
            .O(N__43663),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__9119 (
            .O(N__43658),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__9118 (
            .O(N__43655),
            .I(N__43652));
    LocalMux I__9117 (
            .O(N__43652),
            .I(N__43649));
    Span4Mux_h I__9116 (
            .O(N__43649),
            .I(N__43645));
    InMux I__9115 (
            .O(N__43648),
            .I(N__43642));
    Odrv4 I__9114 (
            .O(N__43645),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__9113 (
            .O(N__43642),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__9112 (
            .O(N__43637),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__9111 (
            .O(N__43634),
            .I(N__43631));
    LocalMux I__9110 (
            .O(N__43631),
            .I(N__43628));
    Span4Mux_h I__9109 (
            .O(N__43628),
            .I(N__43624));
    InMux I__9108 (
            .O(N__43627),
            .I(N__43621));
    Odrv4 I__9107 (
            .O(N__43624),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    LocalMux I__9106 (
            .O(N__43621),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__9105 (
            .O(N__43616),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__9104 (
            .O(N__43613),
            .I(N__43609));
    InMux I__9103 (
            .O(N__43612),
            .I(N__43606));
    InMux I__9102 (
            .O(N__43609),
            .I(N__43603));
    LocalMux I__9101 (
            .O(N__43606),
            .I(N__43600));
    LocalMux I__9100 (
            .O(N__43603),
            .I(N__43597));
    Span4Mux_h I__9099 (
            .O(N__43600),
            .I(N__43594));
    Span4Mux_h I__9098 (
            .O(N__43597),
            .I(N__43591));
    Odrv4 I__9097 (
            .O(N__43594),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__9096 (
            .O(N__43591),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__9095 (
            .O(N__43586),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__9094 (
            .O(N__43583),
            .I(N__43579));
    InMux I__9093 (
            .O(N__43582),
            .I(N__43576));
    LocalMux I__9092 (
            .O(N__43579),
            .I(N__43573));
    LocalMux I__9091 (
            .O(N__43576),
            .I(N__43570));
    Span4Mux_h I__9090 (
            .O(N__43573),
            .I(N__43567));
    Span4Mux_h I__9089 (
            .O(N__43570),
            .I(N__43564));
    Odrv4 I__9088 (
            .O(N__43567),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__9087 (
            .O(N__43564),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__9086 (
            .O(N__43559),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__9085 (
            .O(N__43556),
            .I(N__43553));
    LocalMux I__9084 (
            .O(N__43553),
            .I(N__43549));
    CascadeMux I__9083 (
            .O(N__43552),
            .I(N__43546));
    Span4Mux_v I__9082 (
            .O(N__43549),
            .I(N__43543));
    InMux I__9081 (
            .O(N__43546),
            .I(N__43540));
    Span4Mux_h I__9080 (
            .O(N__43543),
            .I(N__43537));
    LocalMux I__9079 (
            .O(N__43540),
            .I(N__43534));
    Odrv4 I__9078 (
            .O(N__43537),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__9077 (
            .O(N__43534),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__9076 (
            .O(N__43529),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__9075 (
            .O(N__43526),
            .I(N__43523));
    LocalMux I__9074 (
            .O(N__43523),
            .I(N__43520));
    Span4Mux_s1_h I__9073 (
            .O(N__43520),
            .I(N__43516));
    InMux I__9072 (
            .O(N__43519),
            .I(N__43513));
    Span4Mux_h I__9071 (
            .O(N__43516),
            .I(N__43510));
    LocalMux I__9070 (
            .O(N__43513),
            .I(N__43505));
    Span4Mux_h I__9069 (
            .O(N__43510),
            .I(N__43505));
    Odrv4 I__9068 (
            .O(N__43505),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__9067 (
            .O(N__43502),
            .I(N__43499));
    LocalMux I__9066 (
            .O(N__43499),
            .I(N__43496));
    Sp12to4 I__9065 (
            .O(N__43496),
            .I(N__43492));
    InMux I__9064 (
            .O(N__43495),
            .I(N__43489));
    Span12Mux_v I__9063 (
            .O(N__43492),
            .I(N__43486));
    LocalMux I__9062 (
            .O(N__43489),
            .I(N__43483));
    Span12Mux_h I__9061 (
            .O(N__43486),
            .I(N__43480));
    Odrv4 I__9060 (
            .O(N__43483),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    Odrv12 I__9059 (
            .O(N__43480),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    InMux I__9058 (
            .O(N__43475),
            .I(N__43472));
    LocalMux I__9057 (
            .O(N__43472),
            .I(N__43469));
    Span4Mux_v I__9056 (
            .O(N__43469),
            .I(N__43466));
    Span4Mux_v I__9055 (
            .O(N__43466),
            .I(N__43463));
    Span4Mux_v I__9054 (
            .O(N__43463),
            .I(N__43459));
    InMux I__9053 (
            .O(N__43462),
            .I(N__43456));
    Sp12to4 I__9052 (
            .O(N__43459),
            .I(N__43453));
    LocalMux I__9051 (
            .O(N__43456),
            .I(N__43450));
    Span12Mux_s9_h I__9050 (
            .O(N__43453),
            .I(N__43447));
    Odrv4 I__9049 (
            .O(N__43450),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    Odrv12 I__9048 (
            .O(N__43447),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__9047 (
            .O(N__43442),
            .I(N__43439));
    LocalMux I__9046 (
            .O(N__43439),
            .I(N__43436));
    Span12Mux_v I__9045 (
            .O(N__43436),
            .I(N__43432));
    InMux I__9044 (
            .O(N__43435),
            .I(N__43429));
    Span12Mux_h I__9043 (
            .O(N__43432),
            .I(N__43426));
    LocalMux I__9042 (
            .O(N__43429),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    Odrv12 I__9041 (
            .O(N__43426),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__9040 (
            .O(N__43421),
            .I(N__43418));
    LocalMux I__9039 (
            .O(N__43418),
            .I(N__43415));
    Span4Mux_s2_h I__9038 (
            .O(N__43415),
            .I(N__43412));
    Span4Mux_h I__9037 (
            .O(N__43412),
            .I(N__43408));
    InMux I__9036 (
            .O(N__43411),
            .I(N__43405));
    Span4Mux_v I__9035 (
            .O(N__43408),
            .I(N__43402));
    LocalMux I__9034 (
            .O(N__43405),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__9033 (
            .O(N__43402),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__9032 (
            .O(N__43397),
            .I(N__43394));
    LocalMux I__9031 (
            .O(N__43394),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ));
    InMux I__9030 (
            .O(N__43391),
            .I(N__43388));
    LocalMux I__9029 (
            .O(N__43388),
            .I(N__43385));
    Span4Mux_s2_h I__9028 (
            .O(N__43385),
            .I(N__43382));
    Sp12to4 I__9027 (
            .O(N__43382),
            .I(N__43378));
    InMux I__9026 (
            .O(N__43381),
            .I(N__43375));
    Span12Mux_h I__9025 (
            .O(N__43378),
            .I(N__43372));
    LocalMux I__9024 (
            .O(N__43375),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    Odrv12 I__9023 (
            .O(N__43372),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__9022 (
            .O(N__43367),
            .I(N__43364));
    LocalMux I__9021 (
            .O(N__43364),
            .I(N__43361));
    Span12Mux_s7_h I__9020 (
            .O(N__43361),
            .I(N__43357));
    InMux I__9019 (
            .O(N__43360),
            .I(N__43354));
    Span12Mux_v I__9018 (
            .O(N__43357),
            .I(N__43351));
    LocalMux I__9017 (
            .O(N__43354),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    Odrv12 I__9016 (
            .O(N__43351),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    InMux I__9015 (
            .O(N__43346),
            .I(N__43343));
    LocalMux I__9014 (
            .O(N__43343),
            .I(N__43340));
    Span12Mux_v I__9013 (
            .O(N__43340),
            .I(N__43336));
    InMux I__9012 (
            .O(N__43339),
            .I(N__43333));
    Span12Mux_h I__9011 (
            .O(N__43336),
            .I(N__43330));
    LocalMux I__9010 (
            .O(N__43333),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    Odrv12 I__9009 (
            .O(N__43330),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__9008 (
            .O(N__43325),
            .I(N__43322));
    LocalMux I__9007 (
            .O(N__43322),
            .I(N__43319));
    Span4Mux_v I__9006 (
            .O(N__43319),
            .I(N__43316));
    Span4Mux_v I__9005 (
            .O(N__43316),
            .I(N__43313));
    Sp12to4 I__9004 (
            .O(N__43313),
            .I(N__43310));
    Span12Mux_s3_h I__9003 (
            .O(N__43310),
            .I(N__43306));
    InMux I__9002 (
            .O(N__43309),
            .I(N__43303));
    Span12Mux_h I__9001 (
            .O(N__43306),
            .I(N__43300));
    LocalMux I__9000 (
            .O(N__43303),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv12 I__8999 (
            .O(N__43300),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__8998 (
            .O(N__43295),
            .I(N__43292));
    LocalMux I__8997 (
            .O(N__43292),
            .I(N__43289));
    Span4Mux_v I__8996 (
            .O(N__43289),
            .I(N__43286));
    Odrv4 I__8995 (
            .O(N__43286),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__8994 (
            .O(N__43283),
            .I(N__43280));
    LocalMux I__8993 (
            .O(N__43280),
            .I(N__43277));
    Odrv12 I__8992 (
            .O(N__43277),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__8991 (
            .O(N__43274),
            .I(N__43271));
    LocalMux I__8990 (
            .O(N__43271),
            .I(N__43268));
    Span4Mux_v I__8989 (
            .O(N__43268),
            .I(N__43265));
    Odrv4 I__8988 (
            .O(N__43265),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__8987 (
            .O(N__43262),
            .I(N__43259));
    LocalMux I__8986 (
            .O(N__43259),
            .I(N__43256));
    Odrv12 I__8985 (
            .O(N__43256),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__8984 (
            .O(N__43253),
            .I(N__43250));
    LocalMux I__8983 (
            .O(N__43250),
            .I(N__43247));
    Odrv12 I__8982 (
            .O(N__43247),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__8981 (
            .O(N__43244),
            .I(N__43241));
    LocalMux I__8980 (
            .O(N__43241),
            .I(N__43238));
    Odrv12 I__8979 (
            .O(N__43238),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__8978 (
            .O(N__43235),
            .I(N__43232));
    LocalMux I__8977 (
            .O(N__43232),
            .I(N__43229));
    Span4Mux_v I__8976 (
            .O(N__43229),
            .I(N__43226));
    Odrv4 I__8975 (
            .O(N__43226),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__8974 (
            .O(N__43223),
            .I(N__43220));
    LocalMux I__8973 (
            .O(N__43220),
            .I(N__43217));
    Span4Mux_v I__8972 (
            .O(N__43217),
            .I(N__43214));
    Odrv4 I__8971 (
            .O(N__43214),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    CascadeMux I__8970 (
            .O(N__43211),
            .I(N__43208));
    InMux I__8969 (
            .O(N__43208),
            .I(N__43205));
    LocalMux I__8968 (
            .O(N__43205),
            .I(N__43202));
    Odrv12 I__8967 (
            .O(N__43202),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__8966 (
            .O(N__43199),
            .I(N__43196));
    LocalMux I__8965 (
            .O(N__43196),
            .I(N__43193));
    Span4Mux_v I__8964 (
            .O(N__43193),
            .I(N__43190));
    Odrv4 I__8963 (
            .O(N__43190),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__8962 (
            .O(N__43187),
            .I(N__43184));
    LocalMux I__8961 (
            .O(N__43184),
            .I(N__43181));
    Odrv12 I__8960 (
            .O(N__43181),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__8959 (
            .O(N__43178),
            .I(N__43175));
    LocalMux I__8958 (
            .O(N__43175),
            .I(N__43172));
    Span12Mux_v I__8957 (
            .O(N__43172),
            .I(N__43169));
    Odrv12 I__8956 (
            .O(N__43169),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__8955 (
            .O(N__43166),
            .I(N__43163));
    LocalMux I__8954 (
            .O(N__43163),
            .I(N__43160));
    Odrv12 I__8953 (
            .O(N__43160),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__8952 (
            .O(N__43157),
            .I(N__43154));
    LocalMux I__8951 (
            .O(N__43154),
            .I(N__43151));
    Odrv12 I__8950 (
            .O(N__43151),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__8949 (
            .O(N__43148),
            .I(N__43145));
    LocalMux I__8948 (
            .O(N__43145),
            .I(N__43142));
    Odrv12 I__8947 (
            .O(N__43142),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__8946 (
            .O(N__43139),
            .I(N__43136));
    LocalMux I__8945 (
            .O(N__43136),
            .I(N__43133));
    Span4Mux_v I__8944 (
            .O(N__43133),
            .I(N__43130));
    Odrv4 I__8943 (
            .O(N__43130),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__8942 (
            .O(N__43127),
            .I(N__43124));
    LocalMux I__8941 (
            .O(N__43124),
            .I(N__43121));
    Odrv12 I__8940 (
            .O(N__43121),
            .I(\current_shift_inst.un38_control_input_0_s1_3 ));
    CascadeMux I__8939 (
            .O(N__43118),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    CascadeMux I__8938 (
            .O(N__43115),
            .I(N__43112));
    InMux I__8937 (
            .O(N__43112),
            .I(N__43109));
    LocalMux I__8936 (
            .O(N__43109),
            .I(N__43104));
    InMux I__8935 (
            .O(N__43108),
            .I(N__43101));
    InMux I__8934 (
            .O(N__43107),
            .I(N__43098));
    Span4Mux_v I__8933 (
            .O(N__43104),
            .I(N__43095));
    LocalMux I__8932 (
            .O(N__43101),
            .I(N__43092));
    LocalMux I__8931 (
            .O(N__43098),
            .I(N__43089));
    Span4Mux_v I__8930 (
            .O(N__43095),
            .I(N__43085));
    Sp12to4 I__8929 (
            .O(N__43092),
            .I(N__43082));
    Span4Mux_v I__8928 (
            .O(N__43089),
            .I(N__43079));
    InMux I__8927 (
            .O(N__43088),
            .I(N__43076));
    Odrv4 I__8926 (
            .O(N__43085),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv12 I__8925 (
            .O(N__43082),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__8924 (
            .O(N__43079),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__8923 (
            .O(N__43076),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__8922 (
            .O(N__43067),
            .I(N__43063));
    CascadeMux I__8921 (
            .O(N__43066),
            .I(N__43060));
    LocalMux I__8920 (
            .O(N__43063),
            .I(N__43056));
    InMux I__8919 (
            .O(N__43060),
            .I(N__43053));
    InMux I__8918 (
            .O(N__43059),
            .I(N__43050));
    Span4Mux_v I__8917 (
            .O(N__43056),
            .I(N__43047));
    LocalMux I__8916 (
            .O(N__43053),
            .I(N__43044));
    LocalMux I__8915 (
            .O(N__43050),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__8914 (
            .O(N__43047),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__8913 (
            .O(N__43044),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__8912 (
            .O(N__43037),
            .I(N__43034));
    LocalMux I__8911 (
            .O(N__43034),
            .I(N__43031));
    Odrv4 I__8910 (
            .O(N__43031),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__8909 (
            .O(N__43028),
            .I(N__43025));
    LocalMux I__8908 (
            .O(N__43025),
            .I(N__43022));
    Span12Mux_v I__8907 (
            .O(N__43022),
            .I(N__43019));
    Odrv12 I__8906 (
            .O(N__43019),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__8905 (
            .O(N__43016),
            .I(N__43013));
    LocalMux I__8904 (
            .O(N__43013),
            .I(N__43010));
    Odrv12 I__8903 (
            .O(N__43010),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    CascadeMux I__8902 (
            .O(N__43007),
            .I(N__43004));
    InMux I__8901 (
            .O(N__43004),
            .I(N__43001));
    LocalMux I__8900 (
            .O(N__43001),
            .I(N__42998));
    Span4Mux_v I__8899 (
            .O(N__42998),
            .I(N__42995));
    Odrv4 I__8898 (
            .O(N__42995),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    CascadeMux I__8897 (
            .O(N__42992),
            .I(N__42988));
    InMux I__8896 (
            .O(N__42991),
            .I(N__42984));
    InMux I__8895 (
            .O(N__42988),
            .I(N__42981));
    InMux I__8894 (
            .O(N__42987),
            .I(N__42978));
    LocalMux I__8893 (
            .O(N__42984),
            .I(N__42975));
    LocalMux I__8892 (
            .O(N__42981),
            .I(N__42972));
    LocalMux I__8891 (
            .O(N__42978),
            .I(N__42969));
    Span4Mux_v I__8890 (
            .O(N__42975),
            .I(N__42965));
    Span4Mux_v I__8889 (
            .O(N__42972),
            .I(N__42962));
    Span4Mux_v I__8888 (
            .O(N__42969),
            .I(N__42959));
    InMux I__8887 (
            .O(N__42968),
            .I(N__42956));
    Odrv4 I__8886 (
            .O(N__42965),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__8885 (
            .O(N__42962),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__8884 (
            .O(N__42959),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__8883 (
            .O(N__42956),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__8882 (
            .O(N__42947),
            .I(N__42944));
    LocalMux I__8881 (
            .O(N__42944),
            .I(N__42939));
    InMux I__8880 (
            .O(N__42943),
            .I(N__42936));
    InMux I__8879 (
            .O(N__42942),
            .I(N__42933));
    Span4Mux_h I__8878 (
            .O(N__42939),
            .I(N__42930));
    LocalMux I__8877 (
            .O(N__42936),
            .I(N__42927));
    LocalMux I__8876 (
            .O(N__42933),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv4 I__8875 (
            .O(N__42930),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv12 I__8874 (
            .O(N__42927),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__8873 (
            .O(N__42920),
            .I(N__42917));
    LocalMux I__8872 (
            .O(N__42917),
            .I(N__42914));
    Span4Mux_v I__8871 (
            .O(N__42914),
            .I(N__42911));
    Odrv4 I__8870 (
            .O(N__42911),
            .I(\current_shift_inst.un38_control_input_0_s1_4 ));
    InMux I__8869 (
            .O(N__42908),
            .I(N__42905));
    LocalMux I__8868 (
            .O(N__42905),
            .I(N__42902));
    Span4Mux_v I__8867 (
            .O(N__42902),
            .I(N__42899));
    Odrv4 I__8866 (
            .O(N__42899),
            .I(\current_shift_inst.un38_control_input_0_s1_5 ));
    InMux I__8865 (
            .O(N__42896),
            .I(N__42893));
    LocalMux I__8864 (
            .O(N__42893),
            .I(N__42890));
    Odrv12 I__8863 (
            .O(N__42890),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    CascadeMux I__8862 (
            .O(N__42887),
            .I(N__42884));
    InMux I__8861 (
            .O(N__42884),
            .I(N__42881));
    LocalMux I__8860 (
            .O(N__42881),
            .I(N__42877));
    CascadeMux I__8859 (
            .O(N__42880),
            .I(N__42873));
    Span4Mux_v I__8858 (
            .O(N__42877),
            .I(N__42870));
    InMux I__8857 (
            .O(N__42876),
            .I(N__42867));
    InMux I__8856 (
            .O(N__42873),
            .I(N__42864));
    Span4Mux_h I__8855 (
            .O(N__42870),
            .I(N__42861));
    LocalMux I__8854 (
            .O(N__42867),
            .I(N__42858));
    LocalMux I__8853 (
            .O(N__42864),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__8852 (
            .O(N__42861),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv12 I__8851 (
            .O(N__42858),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__8850 (
            .O(N__42851),
            .I(N__42847));
    CascadeMux I__8849 (
            .O(N__42850),
            .I(N__42844));
    LocalMux I__8848 (
            .O(N__42847),
            .I(N__42840));
    InMux I__8847 (
            .O(N__42844),
            .I(N__42837));
    InMux I__8846 (
            .O(N__42843),
            .I(N__42834));
    Span4Mux_h I__8845 (
            .O(N__42840),
            .I(N__42829));
    LocalMux I__8844 (
            .O(N__42837),
            .I(N__42829));
    LocalMux I__8843 (
            .O(N__42834),
            .I(N__42825));
    Span4Mux_v I__8842 (
            .O(N__42829),
            .I(N__42822));
    InMux I__8841 (
            .O(N__42828),
            .I(N__42819));
    Odrv12 I__8840 (
            .O(N__42825),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__8839 (
            .O(N__42822),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__8838 (
            .O(N__42819),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    CascadeMux I__8837 (
            .O(N__42812),
            .I(N__42809));
    InMux I__8836 (
            .O(N__42809),
            .I(N__42806));
    LocalMux I__8835 (
            .O(N__42806),
            .I(N__42803));
    Odrv4 I__8834 (
            .O(N__42803),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    InMux I__8833 (
            .O(N__42800),
            .I(N__42797));
    LocalMux I__8832 (
            .O(N__42797),
            .I(N__42793));
    InMux I__8831 (
            .O(N__42796),
            .I(N__42790));
    Span4Mux_v I__8830 (
            .O(N__42793),
            .I(N__42787));
    LocalMux I__8829 (
            .O(N__42790),
            .I(N__42784));
    Odrv4 I__8828 (
            .O(N__42787),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv12 I__8827 (
            .O(N__42784),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__8826 (
            .O(N__42779),
            .I(N__42758));
    CascadeMux I__8825 (
            .O(N__42778),
            .I(N__42755));
    CascadeMux I__8824 (
            .O(N__42777),
            .I(N__42752));
    CascadeMux I__8823 (
            .O(N__42776),
            .I(N__42749));
    CascadeMux I__8822 (
            .O(N__42775),
            .I(N__42746));
    CascadeMux I__8821 (
            .O(N__42774),
            .I(N__42743));
    CascadeMux I__8820 (
            .O(N__42773),
            .I(N__42740));
    CascadeMux I__8819 (
            .O(N__42772),
            .I(N__42737));
    CascadeMux I__8818 (
            .O(N__42771),
            .I(N__42734));
    CascadeMux I__8817 (
            .O(N__42770),
            .I(N__42731));
    CascadeMux I__8816 (
            .O(N__42769),
            .I(N__42728));
    CascadeMux I__8815 (
            .O(N__42768),
            .I(N__42725));
    CascadeMux I__8814 (
            .O(N__42767),
            .I(N__42722));
    CascadeMux I__8813 (
            .O(N__42766),
            .I(N__42719));
    CascadeMux I__8812 (
            .O(N__42765),
            .I(N__42716));
    CascadeMux I__8811 (
            .O(N__42764),
            .I(N__42713));
    InMux I__8810 (
            .O(N__42763),
            .I(N__42698));
    InMux I__8809 (
            .O(N__42762),
            .I(N__42698));
    InMux I__8808 (
            .O(N__42761),
            .I(N__42695));
    LocalMux I__8807 (
            .O(N__42758),
            .I(N__42692));
    InMux I__8806 (
            .O(N__42755),
            .I(N__42685));
    InMux I__8805 (
            .O(N__42752),
            .I(N__42685));
    InMux I__8804 (
            .O(N__42749),
            .I(N__42685));
    InMux I__8803 (
            .O(N__42746),
            .I(N__42676));
    InMux I__8802 (
            .O(N__42743),
            .I(N__42676));
    InMux I__8801 (
            .O(N__42740),
            .I(N__42676));
    InMux I__8800 (
            .O(N__42737),
            .I(N__42676));
    InMux I__8799 (
            .O(N__42734),
            .I(N__42667));
    InMux I__8798 (
            .O(N__42731),
            .I(N__42667));
    InMux I__8797 (
            .O(N__42728),
            .I(N__42667));
    InMux I__8796 (
            .O(N__42725),
            .I(N__42667));
    InMux I__8795 (
            .O(N__42722),
            .I(N__42658));
    InMux I__8794 (
            .O(N__42719),
            .I(N__42658));
    InMux I__8793 (
            .O(N__42716),
            .I(N__42658));
    InMux I__8792 (
            .O(N__42713),
            .I(N__42658));
    CascadeMux I__8791 (
            .O(N__42712),
            .I(N__42655));
    CascadeMux I__8790 (
            .O(N__42711),
            .I(N__42652));
    CascadeMux I__8789 (
            .O(N__42710),
            .I(N__42649));
    CascadeMux I__8788 (
            .O(N__42709),
            .I(N__42646));
    CascadeMux I__8787 (
            .O(N__42708),
            .I(N__42643));
    CascadeMux I__8786 (
            .O(N__42707),
            .I(N__42640));
    CascadeMux I__8785 (
            .O(N__42706),
            .I(N__42637));
    CascadeMux I__8784 (
            .O(N__42705),
            .I(N__42634));
    InMux I__8783 (
            .O(N__42704),
            .I(N__42627));
    CascadeMux I__8782 (
            .O(N__42703),
            .I(N__42624));
    LocalMux I__8781 (
            .O(N__42698),
            .I(N__42608));
    LocalMux I__8780 (
            .O(N__42695),
            .I(N__42608));
    Span4Mux_s1_h I__8779 (
            .O(N__42692),
            .I(N__42602));
    LocalMux I__8778 (
            .O(N__42685),
            .I(N__42586));
    LocalMux I__8777 (
            .O(N__42676),
            .I(N__42586));
    LocalMux I__8776 (
            .O(N__42667),
            .I(N__42586));
    LocalMux I__8775 (
            .O(N__42658),
            .I(N__42586));
    InMux I__8774 (
            .O(N__42655),
            .I(N__42577));
    InMux I__8773 (
            .O(N__42652),
            .I(N__42577));
    InMux I__8772 (
            .O(N__42649),
            .I(N__42577));
    InMux I__8771 (
            .O(N__42646),
            .I(N__42577));
    InMux I__8770 (
            .O(N__42643),
            .I(N__42568));
    InMux I__8769 (
            .O(N__42640),
            .I(N__42568));
    InMux I__8768 (
            .O(N__42637),
            .I(N__42568));
    InMux I__8767 (
            .O(N__42634),
            .I(N__42568));
    CascadeMux I__8766 (
            .O(N__42633),
            .I(N__42565));
    CascadeMux I__8765 (
            .O(N__42632),
            .I(N__42562));
    CascadeMux I__8764 (
            .O(N__42631),
            .I(N__42559));
    CascadeMux I__8763 (
            .O(N__42630),
            .I(N__42556));
    LocalMux I__8762 (
            .O(N__42627),
            .I(N__42553));
    InMux I__8761 (
            .O(N__42624),
            .I(N__42546));
    CascadeMux I__8760 (
            .O(N__42623),
            .I(N__42543));
    CascadeMux I__8759 (
            .O(N__42622),
            .I(N__42539));
    CascadeMux I__8758 (
            .O(N__42621),
            .I(N__42535));
    CascadeMux I__8757 (
            .O(N__42620),
            .I(N__42531));
    CascadeMux I__8756 (
            .O(N__42619),
            .I(N__42527));
    CascadeMux I__8755 (
            .O(N__42618),
            .I(N__42523));
    CascadeMux I__8754 (
            .O(N__42617),
            .I(N__42519));
    CascadeMux I__8753 (
            .O(N__42616),
            .I(N__42515));
    CascadeMux I__8752 (
            .O(N__42615),
            .I(N__42510));
    CascadeMux I__8751 (
            .O(N__42614),
            .I(N__42506));
    CascadeMux I__8750 (
            .O(N__42613),
            .I(N__42502));
    Span4Mux_s2_h I__8749 (
            .O(N__42608),
            .I(N__42498));
    InMux I__8748 (
            .O(N__42607),
            .I(N__42493));
    InMux I__8747 (
            .O(N__42606),
            .I(N__42493));
    InMux I__8746 (
            .O(N__42605),
            .I(N__42490));
    Span4Mux_h I__8745 (
            .O(N__42602),
            .I(N__42477));
    CascadeMux I__8744 (
            .O(N__42601),
            .I(N__42474));
    CascadeMux I__8743 (
            .O(N__42600),
            .I(N__42471));
    CascadeMux I__8742 (
            .O(N__42599),
            .I(N__42468));
    CascadeMux I__8741 (
            .O(N__42598),
            .I(N__42465));
    CascadeMux I__8740 (
            .O(N__42597),
            .I(N__42462));
    CascadeMux I__8739 (
            .O(N__42596),
            .I(N__42459));
    CascadeMux I__8738 (
            .O(N__42595),
            .I(N__42456));
    Span4Mux_v I__8737 (
            .O(N__42586),
            .I(N__42445));
    LocalMux I__8736 (
            .O(N__42577),
            .I(N__42445));
    LocalMux I__8735 (
            .O(N__42568),
            .I(N__42445));
    InMux I__8734 (
            .O(N__42565),
            .I(N__42440));
    InMux I__8733 (
            .O(N__42562),
            .I(N__42440));
    InMux I__8732 (
            .O(N__42559),
            .I(N__42435));
    InMux I__8731 (
            .O(N__42556),
            .I(N__42435));
    Span4Mux_s1_h I__8730 (
            .O(N__42553),
            .I(N__42432));
    InMux I__8729 (
            .O(N__42552),
            .I(N__42429));
    CascadeMux I__8728 (
            .O(N__42551),
            .I(N__42425));
    CascadeMux I__8727 (
            .O(N__42550),
            .I(N__42421));
    CascadeMux I__8726 (
            .O(N__42549),
            .I(N__42417));
    LocalMux I__8725 (
            .O(N__42546),
            .I(N__42413));
    InMux I__8724 (
            .O(N__42543),
            .I(N__42396));
    InMux I__8723 (
            .O(N__42542),
            .I(N__42396));
    InMux I__8722 (
            .O(N__42539),
            .I(N__42396));
    InMux I__8721 (
            .O(N__42538),
            .I(N__42396));
    InMux I__8720 (
            .O(N__42535),
            .I(N__42396));
    InMux I__8719 (
            .O(N__42534),
            .I(N__42396));
    InMux I__8718 (
            .O(N__42531),
            .I(N__42396));
    InMux I__8717 (
            .O(N__42530),
            .I(N__42396));
    InMux I__8716 (
            .O(N__42527),
            .I(N__42379));
    InMux I__8715 (
            .O(N__42526),
            .I(N__42379));
    InMux I__8714 (
            .O(N__42523),
            .I(N__42379));
    InMux I__8713 (
            .O(N__42522),
            .I(N__42379));
    InMux I__8712 (
            .O(N__42519),
            .I(N__42379));
    InMux I__8711 (
            .O(N__42518),
            .I(N__42379));
    InMux I__8710 (
            .O(N__42515),
            .I(N__42379));
    InMux I__8709 (
            .O(N__42514),
            .I(N__42379));
    InMux I__8708 (
            .O(N__42513),
            .I(N__42364));
    InMux I__8707 (
            .O(N__42510),
            .I(N__42364));
    InMux I__8706 (
            .O(N__42509),
            .I(N__42364));
    InMux I__8705 (
            .O(N__42506),
            .I(N__42364));
    InMux I__8704 (
            .O(N__42505),
            .I(N__42364));
    InMux I__8703 (
            .O(N__42502),
            .I(N__42364));
    InMux I__8702 (
            .O(N__42501),
            .I(N__42364));
    Span4Mux_v I__8701 (
            .O(N__42498),
            .I(N__42353));
    LocalMux I__8700 (
            .O(N__42493),
            .I(N__42348));
    LocalMux I__8699 (
            .O(N__42490),
            .I(N__42348));
    InMux I__8698 (
            .O(N__42489),
            .I(N__42339));
    InMux I__8697 (
            .O(N__42488),
            .I(N__42330));
    InMux I__8696 (
            .O(N__42487),
            .I(N__42330));
    InMux I__8695 (
            .O(N__42486),
            .I(N__42330));
    InMux I__8694 (
            .O(N__42485),
            .I(N__42330));
    InMux I__8693 (
            .O(N__42484),
            .I(N__42319));
    InMux I__8692 (
            .O(N__42483),
            .I(N__42319));
    InMux I__8691 (
            .O(N__42482),
            .I(N__42319));
    InMux I__8690 (
            .O(N__42481),
            .I(N__42319));
    InMux I__8689 (
            .O(N__42480),
            .I(N__42319));
    Span4Mux_h I__8688 (
            .O(N__42477),
            .I(N__42316));
    InMux I__8687 (
            .O(N__42474),
            .I(N__42309));
    InMux I__8686 (
            .O(N__42471),
            .I(N__42309));
    InMux I__8685 (
            .O(N__42468),
            .I(N__42309));
    InMux I__8684 (
            .O(N__42465),
            .I(N__42300));
    InMux I__8683 (
            .O(N__42462),
            .I(N__42300));
    InMux I__8682 (
            .O(N__42459),
            .I(N__42300));
    InMux I__8681 (
            .O(N__42456),
            .I(N__42300));
    CascadeMux I__8680 (
            .O(N__42455),
            .I(N__42297));
    CascadeMux I__8679 (
            .O(N__42454),
            .I(N__42294));
    CascadeMux I__8678 (
            .O(N__42453),
            .I(N__42291));
    CascadeMux I__8677 (
            .O(N__42452),
            .I(N__42288));
    Span4Mux_h I__8676 (
            .O(N__42445),
            .I(N__42281));
    LocalMux I__8675 (
            .O(N__42440),
            .I(N__42281));
    LocalMux I__8674 (
            .O(N__42435),
            .I(N__42281));
    Span4Mux_h I__8673 (
            .O(N__42432),
            .I(N__42278));
    LocalMux I__8672 (
            .O(N__42429),
            .I(N__42275));
    InMux I__8671 (
            .O(N__42428),
            .I(N__42260));
    InMux I__8670 (
            .O(N__42425),
            .I(N__42260));
    InMux I__8669 (
            .O(N__42424),
            .I(N__42260));
    InMux I__8668 (
            .O(N__42421),
            .I(N__42260));
    InMux I__8667 (
            .O(N__42420),
            .I(N__42260));
    InMux I__8666 (
            .O(N__42417),
            .I(N__42260));
    InMux I__8665 (
            .O(N__42416),
            .I(N__42260));
    Span4Mux_v I__8664 (
            .O(N__42413),
            .I(N__42251));
    LocalMux I__8663 (
            .O(N__42396),
            .I(N__42251));
    LocalMux I__8662 (
            .O(N__42379),
            .I(N__42251));
    LocalMux I__8661 (
            .O(N__42364),
            .I(N__42251));
    CascadeMux I__8660 (
            .O(N__42363),
            .I(N__42248));
    CascadeMux I__8659 (
            .O(N__42362),
            .I(N__42245));
    CascadeMux I__8658 (
            .O(N__42361),
            .I(N__42242));
    CascadeMux I__8657 (
            .O(N__42360),
            .I(N__42239));
    CascadeMux I__8656 (
            .O(N__42359),
            .I(N__42236));
    CascadeMux I__8655 (
            .O(N__42358),
            .I(N__42233));
    CascadeMux I__8654 (
            .O(N__42357),
            .I(N__42230));
    CascadeMux I__8653 (
            .O(N__42356),
            .I(N__42227));
    Span4Mux_v I__8652 (
            .O(N__42353),
            .I(N__42213));
    Span4Mux_s2_h I__8651 (
            .O(N__42348),
            .I(N__42213));
    InMux I__8650 (
            .O(N__42347),
            .I(N__42206));
    InMux I__8649 (
            .O(N__42346),
            .I(N__42206));
    InMux I__8648 (
            .O(N__42345),
            .I(N__42203));
    CascadeMux I__8647 (
            .O(N__42344),
            .I(N__42199));
    CascadeMux I__8646 (
            .O(N__42343),
            .I(N__42195));
    CascadeMux I__8645 (
            .O(N__42342),
            .I(N__42191));
    LocalMux I__8644 (
            .O(N__42339),
            .I(N__42182));
    LocalMux I__8643 (
            .O(N__42330),
            .I(N__42182));
    LocalMux I__8642 (
            .O(N__42319),
            .I(N__42182));
    Span4Mux_h I__8641 (
            .O(N__42316),
            .I(N__42179));
    LocalMux I__8640 (
            .O(N__42309),
            .I(N__42174));
    LocalMux I__8639 (
            .O(N__42300),
            .I(N__42174));
    InMux I__8638 (
            .O(N__42297),
            .I(N__42165));
    InMux I__8637 (
            .O(N__42294),
            .I(N__42165));
    InMux I__8636 (
            .O(N__42291),
            .I(N__42165));
    InMux I__8635 (
            .O(N__42288),
            .I(N__42165));
    Span4Mux_v I__8634 (
            .O(N__42281),
            .I(N__42162));
    Span4Mux_h I__8633 (
            .O(N__42278),
            .I(N__42153));
    Span4Mux_v I__8632 (
            .O(N__42275),
            .I(N__42153));
    LocalMux I__8631 (
            .O(N__42260),
            .I(N__42153));
    Span4Mux_v I__8630 (
            .O(N__42251),
            .I(N__42153));
    InMux I__8629 (
            .O(N__42248),
            .I(N__42144));
    InMux I__8628 (
            .O(N__42245),
            .I(N__42144));
    InMux I__8627 (
            .O(N__42242),
            .I(N__42144));
    InMux I__8626 (
            .O(N__42239),
            .I(N__42144));
    InMux I__8625 (
            .O(N__42236),
            .I(N__42135));
    InMux I__8624 (
            .O(N__42233),
            .I(N__42135));
    InMux I__8623 (
            .O(N__42230),
            .I(N__42135));
    InMux I__8622 (
            .O(N__42227),
            .I(N__42135));
    CascadeMux I__8621 (
            .O(N__42226),
            .I(N__42132));
    CascadeMux I__8620 (
            .O(N__42225),
            .I(N__42129));
    CascadeMux I__8619 (
            .O(N__42224),
            .I(N__42126));
    CascadeMux I__8618 (
            .O(N__42223),
            .I(N__42123));
    CascadeMux I__8617 (
            .O(N__42222),
            .I(N__42120));
    CascadeMux I__8616 (
            .O(N__42221),
            .I(N__42117));
    CascadeMux I__8615 (
            .O(N__42220),
            .I(N__42114));
    CascadeMux I__8614 (
            .O(N__42219),
            .I(N__42111));
    InMux I__8613 (
            .O(N__42218),
            .I(N__42107));
    Span4Mux_h I__8612 (
            .O(N__42213),
            .I(N__42103));
    InMux I__8611 (
            .O(N__42212),
            .I(N__42100));
    InMux I__8610 (
            .O(N__42211),
            .I(N__42092));
    LocalMux I__8609 (
            .O(N__42206),
            .I(N__42086));
    LocalMux I__8608 (
            .O(N__42203),
            .I(N__42086));
    InMux I__8607 (
            .O(N__42202),
            .I(N__42071));
    InMux I__8606 (
            .O(N__42199),
            .I(N__42071));
    InMux I__8605 (
            .O(N__42198),
            .I(N__42071));
    InMux I__8604 (
            .O(N__42195),
            .I(N__42071));
    InMux I__8603 (
            .O(N__42194),
            .I(N__42071));
    InMux I__8602 (
            .O(N__42191),
            .I(N__42071));
    InMux I__8601 (
            .O(N__42190),
            .I(N__42071));
    CascadeMux I__8600 (
            .O(N__42189),
            .I(N__42068));
    Span4Mux_v I__8599 (
            .O(N__42182),
            .I(N__42065));
    Span4Mux_h I__8598 (
            .O(N__42179),
            .I(N__42062));
    Span4Mux_v I__8597 (
            .O(N__42174),
            .I(N__42057));
    LocalMux I__8596 (
            .O(N__42165),
            .I(N__42057));
    Span4Mux_v I__8595 (
            .O(N__42162),
            .I(N__42048));
    Span4Mux_h I__8594 (
            .O(N__42153),
            .I(N__42048));
    LocalMux I__8593 (
            .O(N__42144),
            .I(N__42048));
    LocalMux I__8592 (
            .O(N__42135),
            .I(N__42048));
    InMux I__8591 (
            .O(N__42132),
            .I(N__42039));
    InMux I__8590 (
            .O(N__42129),
            .I(N__42039));
    InMux I__8589 (
            .O(N__42126),
            .I(N__42039));
    InMux I__8588 (
            .O(N__42123),
            .I(N__42039));
    InMux I__8587 (
            .O(N__42120),
            .I(N__42034));
    InMux I__8586 (
            .O(N__42117),
            .I(N__42034));
    InMux I__8585 (
            .O(N__42114),
            .I(N__42029));
    InMux I__8584 (
            .O(N__42111),
            .I(N__42029));
    InMux I__8583 (
            .O(N__42110),
            .I(N__42026));
    LocalMux I__8582 (
            .O(N__42107),
            .I(N__42023));
    InMux I__8581 (
            .O(N__42106),
            .I(N__42020));
    Span4Mux_h I__8580 (
            .O(N__42103),
            .I(N__42016));
    LocalMux I__8579 (
            .O(N__42100),
            .I(N__42013));
    InMux I__8578 (
            .O(N__42099),
            .I(N__42008));
    InMux I__8577 (
            .O(N__42098),
            .I(N__42008));
    InMux I__8576 (
            .O(N__42097),
            .I(N__42005));
    CascadeMux I__8575 (
            .O(N__42096),
            .I(N__41993));
    CascadeMux I__8574 (
            .O(N__42095),
            .I(N__41990));
    LocalMux I__8573 (
            .O(N__42092),
            .I(N__41986));
    InMux I__8572 (
            .O(N__42091),
            .I(N__41983));
    Span4Mux_s3_h I__8571 (
            .O(N__42086),
            .I(N__41980));
    LocalMux I__8570 (
            .O(N__42071),
            .I(N__41977));
    InMux I__8569 (
            .O(N__42068),
            .I(N__41974));
    Span4Mux_v I__8568 (
            .O(N__42065),
            .I(N__41971));
    Span4Mux_v I__8567 (
            .O(N__42062),
            .I(N__41966));
    Span4Mux_v I__8566 (
            .O(N__42057),
            .I(N__41966));
    Span4Mux_h I__8565 (
            .O(N__42048),
            .I(N__41957));
    LocalMux I__8564 (
            .O(N__42039),
            .I(N__41957));
    LocalMux I__8563 (
            .O(N__42034),
            .I(N__41957));
    LocalMux I__8562 (
            .O(N__42029),
            .I(N__41957));
    LocalMux I__8561 (
            .O(N__42026),
            .I(N__41950));
    Span4Mux_s1_v I__8560 (
            .O(N__42023),
            .I(N__41950));
    LocalMux I__8559 (
            .O(N__42020),
            .I(N__41950));
    InMux I__8558 (
            .O(N__42019),
            .I(N__41947));
    Span4Mux_h I__8557 (
            .O(N__42016),
            .I(N__41944));
    Span4Mux_s3_h I__8556 (
            .O(N__42013),
            .I(N__41941));
    LocalMux I__8555 (
            .O(N__42008),
            .I(N__41936));
    LocalMux I__8554 (
            .O(N__42005),
            .I(N__41936));
    InMux I__8553 (
            .O(N__42004),
            .I(N__41927));
    InMux I__8552 (
            .O(N__42003),
            .I(N__41927));
    InMux I__8551 (
            .O(N__42002),
            .I(N__41927));
    InMux I__8550 (
            .O(N__42001),
            .I(N__41927));
    InMux I__8549 (
            .O(N__42000),
            .I(N__41916));
    InMux I__8548 (
            .O(N__41999),
            .I(N__41916));
    InMux I__8547 (
            .O(N__41998),
            .I(N__41916));
    InMux I__8546 (
            .O(N__41997),
            .I(N__41916));
    InMux I__8545 (
            .O(N__41996),
            .I(N__41916));
    InMux I__8544 (
            .O(N__41993),
            .I(N__41909));
    InMux I__8543 (
            .O(N__41990),
            .I(N__41909));
    InMux I__8542 (
            .O(N__41989),
            .I(N__41909));
    Span12Mux_s10_h I__8541 (
            .O(N__41986),
            .I(N__41906));
    LocalMux I__8540 (
            .O(N__41983),
            .I(N__41903));
    Span4Mux_v I__8539 (
            .O(N__41980),
            .I(N__41896));
    Span4Mux_s3_h I__8538 (
            .O(N__41977),
            .I(N__41896));
    LocalMux I__8537 (
            .O(N__41974),
            .I(N__41896));
    Span4Mux_v I__8536 (
            .O(N__41971),
            .I(N__41893));
    Span4Mux_v I__8535 (
            .O(N__41966),
            .I(N__41888));
    Span4Mux_v I__8534 (
            .O(N__41957),
            .I(N__41888));
    Span4Mux_v I__8533 (
            .O(N__41950),
            .I(N__41883));
    LocalMux I__8532 (
            .O(N__41947),
            .I(N__41883));
    Span4Mux_h I__8531 (
            .O(N__41944),
            .I(N__41880));
    Span4Mux_v I__8530 (
            .O(N__41941),
            .I(N__41875));
    Span4Mux_s3_h I__8529 (
            .O(N__41936),
            .I(N__41875));
    LocalMux I__8528 (
            .O(N__41927),
            .I(N__41870));
    LocalMux I__8527 (
            .O(N__41916),
            .I(N__41870));
    LocalMux I__8526 (
            .O(N__41909),
            .I(N__41867));
    Span12Mux_h I__8525 (
            .O(N__41906),
            .I(N__41864));
    Span4Mux_s3_h I__8524 (
            .O(N__41903),
            .I(N__41861));
    Span4Mux_v I__8523 (
            .O(N__41896),
            .I(N__41858));
    Span4Mux_v I__8522 (
            .O(N__41893),
            .I(N__41851));
    Span4Mux_h I__8521 (
            .O(N__41888),
            .I(N__41851));
    Span4Mux_v I__8520 (
            .O(N__41883),
            .I(N__41851));
    Span4Mux_h I__8519 (
            .O(N__41880),
            .I(N__41842));
    Span4Mux_v I__8518 (
            .O(N__41875),
            .I(N__41842));
    Span4Mux_s3_h I__8517 (
            .O(N__41870),
            .I(N__41842));
    Span4Mux_s3_h I__8516 (
            .O(N__41867),
            .I(N__41842));
    Odrv12 I__8515 (
            .O(N__41864),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8514 (
            .O(N__41861),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8513 (
            .O(N__41858),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8512 (
            .O(N__41851),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8511 (
            .O(N__41842),
            .I(CONSTANT_ONE_NET));
    InMux I__8510 (
            .O(N__41831),
            .I(N__41828));
    LocalMux I__8509 (
            .O(N__41828),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    CascadeMux I__8508 (
            .O(N__41825),
            .I(N__41822));
    InMux I__8507 (
            .O(N__41822),
            .I(N__41817));
    CascadeMux I__8506 (
            .O(N__41821),
            .I(N__41814));
    InMux I__8505 (
            .O(N__41820),
            .I(N__41811));
    LocalMux I__8504 (
            .O(N__41817),
            .I(N__41808));
    InMux I__8503 (
            .O(N__41814),
            .I(N__41805));
    LocalMux I__8502 (
            .O(N__41811),
            .I(N__41802));
    Span4Mux_v I__8501 (
            .O(N__41808),
            .I(N__41798));
    LocalMux I__8500 (
            .O(N__41805),
            .I(N__41795));
    Span4Mux_v I__8499 (
            .O(N__41802),
            .I(N__41792));
    InMux I__8498 (
            .O(N__41801),
            .I(N__41789));
    Odrv4 I__8497 (
            .O(N__41798),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv12 I__8496 (
            .O(N__41795),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__8495 (
            .O(N__41792),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__8494 (
            .O(N__41789),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__8493 (
            .O(N__41780),
            .I(N__41777));
    LocalMux I__8492 (
            .O(N__41777),
            .I(N__41772));
    InMux I__8491 (
            .O(N__41776),
            .I(N__41769));
    InMux I__8490 (
            .O(N__41775),
            .I(N__41766));
    Span12Mux_s11_h I__8489 (
            .O(N__41772),
            .I(N__41763));
    LocalMux I__8488 (
            .O(N__41769),
            .I(N__41760));
    LocalMux I__8487 (
            .O(N__41766),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv12 I__8486 (
            .O(N__41763),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__8485 (
            .O(N__41760),
            .I(\current_shift_inst.un4_control_input1_20 ));
    CascadeMux I__8484 (
            .O(N__41753),
            .I(N__41750));
    InMux I__8483 (
            .O(N__41750),
            .I(N__41746));
    InMux I__8482 (
            .O(N__41749),
            .I(N__41742));
    LocalMux I__8481 (
            .O(N__41746),
            .I(N__41739));
    InMux I__8480 (
            .O(N__41745),
            .I(N__41736));
    LocalMux I__8479 (
            .O(N__41742),
            .I(N__41733));
    Span4Mux_h I__8478 (
            .O(N__41739),
            .I(N__41728));
    LocalMux I__8477 (
            .O(N__41736),
            .I(N__41728));
    Odrv4 I__8476 (
            .O(N__41733),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__8475 (
            .O(N__41728),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__8474 (
            .O(N__41723),
            .I(N__41719));
    CascadeMux I__8473 (
            .O(N__41722),
            .I(N__41715));
    InMux I__8472 (
            .O(N__41719),
            .I(N__41712));
    InMux I__8471 (
            .O(N__41718),
            .I(N__41709));
    InMux I__8470 (
            .O(N__41715),
            .I(N__41706));
    LocalMux I__8469 (
            .O(N__41712),
            .I(N__41703));
    LocalMux I__8468 (
            .O(N__41709),
            .I(N__41700));
    LocalMux I__8467 (
            .O(N__41706),
            .I(N__41697));
    Span4Mux_h I__8466 (
            .O(N__41703),
            .I(N__41691));
    Span4Mux_v I__8465 (
            .O(N__41700),
            .I(N__41691));
    Span4Mux_v I__8464 (
            .O(N__41697),
            .I(N__41688));
    InMux I__8463 (
            .O(N__41696),
            .I(N__41685));
    Odrv4 I__8462 (
            .O(N__41691),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__8461 (
            .O(N__41688),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__8460 (
            .O(N__41685),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    CascadeMux I__8459 (
            .O(N__41678),
            .I(N__41675));
    InMux I__8458 (
            .O(N__41675),
            .I(N__41671));
    InMux I__8457 (
            .O(N__41674),
            .I(N__41667));
    LocalMux I__8456 (
            .O(N__41671),
            .I(N__41664));
    InMux I__8455 (
            .O(N__41670),
            .I(N__41661));
    LocalMux I__8454 (
            .O(N__41667),
            .I(N__41658));
    Span4Mux_v I__8453 (
            .O(N__41664),
            .I(N__41654));
    LocalMux I__8452 (
            .O(N__41661),
            .I(N__41649));
    Sp12to4 I__8451 (
            .O(N__41658),
            .I(N__41649));
    InMux I__8450 (
            .O(N__41657),
            .I(N__41646));
    Odrv4 I__8449 (
            .O(N__41654),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv12 I__8448 (
            .O(N__41649),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__8447 (
            .O(N__41646),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__8446 (
            .O(N__41639),
            .I(N__41635));
    CascadeMux I__8445 (
            .O(N__41638),
            .I(N__41631));
    LocalMux I__8444 (
            .O(N__41635),
            .I(N__41628));
    InMux I__8443 (
            .O(N__41634),
            .I(N__41625));
    InMux I__8442 (
            .O(N__41631),
            .I(N__41622));
    Span4Mux_h I__8441 (
            .O(N__41628),
            .I(N__41619));
    LocalMux I__8440 (
            .O(N__41625),
            .I(N__41616));
    LocalMux I__8439 (
            .O(N__41622),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__8438 (
            .O(N__41619),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv12 I__8437 (
            .O(N__41616),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__8436 (
            .O(N__41609),
            .I(N__41606));
    LocalMux I__8435 (
            .O(N__41606),
            .I(N__41603));
    Odrv4 I__8434 (
            .O(N__41603),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__8433 (
            .O(N__41600),
            .I(N__41597));
    LocalMux I__8432 (
            .O(N__41597),
            .I(N__41594));
    Odrv4 I__8431 (
            .O(N__41594),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    CascadeMux I__8430 (
            .O(N__41591),
            .I(N__41588));
    InMux I__8429 (
            .O(N__41588),
            .I(N__41585));
    LocalMux I__8428 (
            .O(N__41585),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__8427 (
            .O(N__41582),
            .I(bfn_16_16_0_));
    InMux I__8426 (
            .O(N__41579),
            .I(N__41576));
    LocalMux I__8425 (
            .O(N__41576),
            .I(N__41573));
    Span4Mux_h I__8424 (
            .O(N__41573),
            .I(N__41570));
    Odrv4 I__8423 (
            .O(N__41570),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__8422 (
            .O(N__41567),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__8421 (
            .O(N__41564),
            .I(N__41561));
    InMux I__8420 (
            .O(N__41561),
            .I(N__41558));
    LocalMux I__8419 (
            .O(N__41558),
            .I(N__41555));
    Span4Mux_h I__8418 (
            .O(N__41555),
            .I(N__41552));
    Odrv4 I__8417 (
            .O(N__41552),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__8416 (
            .O(N__41549),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__8415 (
            .O(N__41546),
            .I(N__41543));
    LocalMux I__8414 (
            .O(N__41543),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__8413 (
            .O(N__41540),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    CascadeMux I__8412 (
            .O(N__41537),
            .I(N__41534));
    InMux I__8411 (
            .O(N__41534),
            .I(N__41531));
    LocalMux I__8410 (
            .O(N__41531),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__8409 (
            .O(N__41528),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__8408 (
            .O(N__41525),
            .I(N__41522));
    LocalMux I__8407 (
            .O(N__41522),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__8406 (
            .O(N__41519),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    CascadeMux I__8405 (
            .O(N__41516),
            .I(N__41513));
    InMux I__8404 (
            .O(N__41513),
            .I(N__41510));
    LocalMux I__8403 (
            .O(N__41510),
            .I(N__41507));
    Span4Mux_h I__8402 (
            .O(N__41507),
            .I(N__41504));
    Odrv4 I__8401 (
            .O(N__41504),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    InMux I__8400 (
            .O(N__41501),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__8399 (
            .O(N__41498),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__8398 (
            .O(N__41495),
            .I(N__41492));
    LocalMux I__8397 (
            .O(N__41492),
            .I(N__41489));
    Odrv4 I__8396 (
            .O(N__41489),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    CascadeMux I__8395 (
            .O(N__41486),
            .I(N__41483));
    InMux I__8394 (
            .O(N__41483),
            .I(N__41480));
    LocalMux I__8393 (
            .O(N__41480),
            .I(N__41477));
    Span4Mux_h I__8392 (
            .O(N__41477),
            .I(N__41474));
    Odrv4 I__8391 (
            .O(N__41474),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    InMux I__8390 (
            .O(N__41471),
            .I(bfn_16_15_0_));
    InMux I__8389 (
            .O(N__41468),
            .I(N__41465));
    LocalMux I__8388 (
            .O(N__41465),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    InMux I__8387 (
            .O(N__41462),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    CascadeMux I__8386 (
            .O(N__41459),
            .I(N__41456));
    InMux I__8385 (
            .O(N__41456),
            .I(N__41453));
    LocalMux I__8384 (
            .O(N__41453),
            .I(N__41450));
    Odrv4 I__8383 (
            .O(N__41450),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    InMux I__8382 (
            .O(N__41447),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    InMux I__8381 (
            .O(N__41444),
            .I(N__41441));
    LocalMux I__8380 (
            .O(N__41441),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    InMux I__8379 (
            .O(N__41438),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    CascadeMux I__8378 (
            .O(N__41435),
            .I(N__41432));
    InMux I__8377 (
            .O(N__41432),
            .I(N__41429));
    LocalMux I__8376 (
            .O(N__41429),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__8375 (
            .O(N__41426),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__8374 (
            .O(N__41423),
            .I(N__41420));
    LocalMux I__8373 (
            .O(N__41420),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__8372 (
            .O(N__41417),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    CascadeMux I__8371 (
            .O(N__41414),
            .I(N__41411));
    InMux I__8370 (
            .O(N__41411),
            .I(N__41408));
    LocalMux I__8369 (
            .O(N__41408),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__8368 (
            .O(N__41405),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__8367 (
            .O(N__41402),
            .I(N__41399));
    LocalMux I__8366 (
            .O(N__41399),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__8365 (
            .O(N__41396),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__8364 (
            .O(N__41393),
            .I(N__41390));
    LocalMux I__8363 (
            .O(N__41390),
            .I(N__41387));
    Odrv12 I__8362 (
            .O(N__41387),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    InMux I__8361 (
            .O(N__41384),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    CascadeMux I__8360 (
            .O(N__41381),
            .I(N__41378));
    InMux I__8359 (
            .O(N__41378),
            .I(N__41375));
    LocalMux I__8358 (
            .O(N__41375),
            .I(N__41372));
    Span4Mux_h I__8357 (
            .O(N__41372),
            .I(N__41369));
    Span4Mux_v I__8356 (
            .O(N__41369),
            .I(N__41366));
    Odrv4 I__8355 (
            .O(N__41366),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__8354 (
            .O(N__41363),
            .I(bfn_16_14_0_));
    InMux I__8353 (
            .O(N__41360),
            .I(N__41357));
    LocalMux I__8352 (
            .O(N__41357),
            .I(N__41354));
    Span4Mux_h I__8351 (
            .O(N__41354),
            .I(N__41351));
    Odrv4 I__8350 (
            .O(N__41351),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__8349 (
            .O(N__41348),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__8348 (
            .O(N__41345),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__8347 (
            .O(N__41342),
            .I(N__41339));
    LocalMux I__8346 (
            .O(N__41339),
            .I(N__41336));
    Span4Mux_h I__8345 (
            .O(N__41336),
            .I(N__41333));
    Odrv4 I__8344 (
            .O(N__41333),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    InMux I__8343 (
            .O(N__41330),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    CascadeMux I__8342 (
            .O(N__41327),
            .I(N__41324));
    InMux I__8341 (
            .O(N__41324),
            .I(N__41321));
    LocalMux I__8340 (
            .O(N__41321),
            .I(N__41318));
    Span4Mux_h I__8339 (
            .O(N__41318),
            .I(N__41315));
    Odrv4 I__8338 (
            .O(N__41315),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    InMux I__8337 (
            .O(N__41312),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__8336 (
            .O(N__41309),
            .I(N__41306));
    LocalMux I__8335 (
            .O(N__41306),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    InMux I__8334 (
            .O(N__41303),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    CascadeMux I__8333 (
            .O(N__41300),
            .I(N__41297));
    InMux I__8332 (
            .O(N__41297),
            .I(N__41294));
    LocalMux I__8331 (
            .O(N__41294),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    InMux I__8330 (
            .O(N__41291),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__8329 (
            .O(N__41288),
            .I(N__41285));
    LocalMux I__8328 (
            .O(N__41285),
            .I(N__41282));
    Span4Mux_h I__8327 (
            .O(N__41282),
            .I(N__41279));
    Odrv4 I__8326 (
            .O(N__41279),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    InMux I__8325 (
            .O(N__41276),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__8324 (
            .O(N__41273),
            .I(N__41269));
    InMux I__8323 (
            .O(N__41272),
            .I(N__41265));
    LocalMux I__8322 (
            .O(N__41269),
            .I(N__41262));
    InMux I__8321 (
            .O(N__41268),
            .I(N__41259));
    LocalMux I__8320 (
            .O(N__41265),
            .I(N__41256));
    Span4Mux_h I__8319 (
            .O(N__41262),
            .I(N__41252));
    LocalMux I__8318 (
            .O(N__41259),
            .I(N__41247));
    Sp12to4 I__8317 (
            .O(N__41256),
            .I(N__41247));
    InMux I__8316 (
            .O(N__41255),
            .I(N__41244));
    Odrv4 I__8315 (
            .O(N__41252),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv12 I__8314 (
            .O(N__41247),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__8313 (
            .O(N__41244),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__8312 (
            .O(N__41237),
            .I(N__41234));
    LocalMux I__8311 (
            .O(N__41234),
            .I(N__41231));
    Span4Mux_v I__8310 (
            .O(N__41231),
            .I(N__41228));
    Odrv4 I__8309 (
            .O(N__41228),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    CascadeMux I__8308 (
            .O(N__41225),
            .I(N__41222));
    InMux I__8307 (
            .O(N__41222),
            .I(N__41219));
    LocalMux I__8306 (
            .O(N__41219),
            .I(N__41216));
    Span4Mux_h I__8305 (
            .O(N__41216),
            .I(N__41213));
    Span4Mux_h I__8304 (
            .O(N__41213),
            .I(N__41210));
    Odrv4 I__8303 (
            .O(N__41210),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__8302 (
            .O(N__41207),
            .I(N__41204));
    InMux I__8301 (
            .O(N__41204),
            .I(N__41201));
    LocalMux I__8300 (
            .O(N__41201),
            .I(N__41198));
    Odrv12 I__8299 (
            .O(N__41198),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__8298 (
            .O(N__41195),
            .I(\current_shift_inst.un38_control_input_cry_2_s1 ));
    CascadeMux I__8297 (
            .O(N__41192),
            .I(N__41189));
    InMux I__8296 (
            .O(N__41189),
            .I(N__41186));
    LocalMux I__8295 (
            .O(N__41186),
            .I(N__41183));
    Odrv4 I__8294 (
            .O(N__41183),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ));
    InMux I__8293 (
            .O(N__41180),
            .I(\current_shift_inst.un38_control_input_cry_3_s1 ));
    InMux I__8292 (
            .O(N__41177),
            .I(N__41174));
    LocalMux I__8291 (
            .O(N__41174),
            .I(N__41171));
    Span4Mux_h I__8290 (
            .O(N__41171),
            .I(N__41168));
    Odrv4 I__8289 (
            .O(N__41168),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ));
    InMux I__8288 (
            .O(N__41165),
            .I(\current_shift_inst.un38_control_input_cry_4_s1 ));
    CascadeMux I__8287 (
            .O(N__41162),
            .I(N__41159));
    InMux I__8286 (
            .O(N__41159),
            .I(N__41156));
    LocalMux I__8285 (
            .O(N__41156),
            .I(N__41153));
    Span4Mux_h I__8284 (
            .O(N__41153),
            .I(N__41150));
    Span4Mux_h I__8283 (
            .O(N__41150),
            .I(N__41147));
    Odrv4 I__8282 (
            .O(N__41147),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__8281 (
            .O(N__41144),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__8280 (
            .O(N__41141),
            .I(N__41137));
    InMux I__8279 (
            .O(N__41140),
            .I(N__41134));
    LocalMux I__8278 (
            .O(N__41137),
            .I(N__41128));
    LocalMux I__8277 (
            .O(N__41134),
            .I(N__41128));
    InMux I__8276 (
            .O(N__41133),
            .I(N__41125));
    Span4Mux_h I__8275 (
            .O(N__41128),
            .I(N__41122));
    LocalMux I__8274 (
            .O(N__41125),
            .I(N__41119));
    Span4Mux_v I__8273 (
            .O(N__41122),
            .I(N__41116));
    Span12Mux_h I__8272 (
            .O(N__41119),
            .I(N__41113));
    Span4Mux_v I__8271 (
            .O(N__41116),
            .I(N__41110));
    Odrv12 I__8270 (
            .O(N__41113),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__8269 (
            .O(N__41110),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__8268 (
            .O(N__41105),
            .I(N__41100));
    InMux I__8267 (
            .O(N__41104),
            .I(N__41095));
    InMux I__8266 (
            .O(N__41103),
            .I(N__41095));
    LocalMux I__8265 (
            .O(N__41100),
            .I(N__41089));
    LocalMux I__8264 (
            .O(N__41095),
            .I(N__41089));
    InMux I__8263 (
            .O(N__41094),
            .I(N__41086));
    Span12Mux_s11_h I__8262 (
            .O(N__41089),
            .I(N__41083));
    LocalMux I__8261 (
            .O(N__41086),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__8260 (
            .O(N__41083),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__8259 (
            .O(N__41078),
            .I(N__41075));
    LocalMux I__8258 (
            .O(N__41075),
            .I(N__41069));
    InMux I__8257 (
            .O(N__41074),
            .I(N__41066));
    InMux I__8256 (
            .O(N__41073),
            .I(N__41063));
    InMux I__8255 (
            .O(N__41072),
            .I(N__41060));
    Span4Mux_v I__8254 (
            .O(N__41069),
            .I(N__41057));
    LocalMux I__8253 (
            .O(N__41066),
            .I(N__41054));
    LocalMux I__8252 (
            .O(N__41063),
            .I(N__41050));
    LocalMux I__8251 (
            .O(N__41060),
            .I(N__41047));
    Sp12to4 I__8250 (
            .O(N__41057),
            .I(N__41044));
    Span4Mux_v I__8249 (
            .O(N__41054),
            .I(N__41041));
    InMux I__8248 (
            .O(N__41053),
            .I(N__41038));
    Span4Mux_v I__8247 (
            .O(N__41050),
            .I(N__41035));
    Span4Mux_h I__8246 (
            .O(N__41047),
            .I(N__41032));
    Odrv12 I__8245 (
            .O(N__41044),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__8244 (
            .O(N__41041),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__8243 (
            .O(N__41038),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__8242 (
            .O(N__41035),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__8241 (
            .O(N__41032),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__8240 (
            .O(N__41021),
            .I(N__41017));
    InMux I__8239 (
            .O(N__41020),
            .I(N__41013));
    LocalMux I__8238 (
            .O(N__41017),
            .I(N__41010));
    CascadeMux I__8237 (
            .O(N__41016),
            .I(N__41007));
    LocalMux I__8236 (
            .O(N__41013),
            .I(N__41004));
    Span4Mux_v I__8235 (
            .O(N__41010),
            .I(N__41001));
    InMux I__8234 (
            .O(N__41007),
            .I(N__40998));
    Span4Mux_v I__8233 (
            .O(N__41004),
            .I(N__40993));
    Span4Mux_h I__8232 (
            .O(N__41001),
            .I(N__40993));
    LocalMux I__8231 (
            .O(N__40998),
            .I(N__40990));
    Odrv4 I__8230 (
            .O(N__40993),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ));
    Odrv4 I__8229 (
            .O(N__40990),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ));
    InMux I__8228 (
            .O(N__40985),
            .I(N__40982));
    LocalMux I__8227 (
            .O(N__40982),
            .I(N__40979));
    Span4Mux_h I__8226 (
            .O(N__40979),
            .I(N__40976));
    Span4Mux_h I__8225 (
            .O(N__40976),
            .I(N__40973));
    Span4Mux_v I__8224 (
            .O(N__40973),
            .I(N__40970));
    Odrv4 I__8223 (
            .O(N__40970),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ));
    CEMux I__8222 (
            .O(N__40967),
            .I(N__40963));
    CEMux I__8221 (
            .O(N__40966),
            .I(N__40960));
    LocalMux I__8220 (
            .O(N__40963),
            .I(N__40957));
    LocalMux I__8219 (
            .O(N__40960),
            .I(N__40951));
    Span4Mux_v I__8218 (
            .O(N__40957),
            .I(N__40948));
    CEMux I__8217 (
            .O(N__40956),
            .I(N__40945));
    CEMux I__8216 (
            .O(N__40955),
            .I(N__40942));
    CEMux I__8215 (
            .O(N__40954),
            .I(N__40938));
    Span4Mux_h I__8214 (
            .O(N__40951),
            .I(N__40934));
    Span4Mux_v I__8213 (
            .O(N__40948),
            .I(N__40931));
    LocalMux I__8212 (
            .O(N__40945),
            .I(N__40928));
    LocalMux I__8211 (
            .O(N__40942),
            .I(N__40925));
    CEMux I__8210 (
            .O(N__40941),
            .I(N__40922));
    LocalMux I__8209 (
            .O(N__40938),
            .I(N__40919));
    CEMux I__8208 (
            .O(N__40937),
            .I(N__40916));
    Span4Mux_v I__8207 (
            .O(N__40934),
            .I(N__40912));
    Span4Mux_h I__8206 (
            .O(N__40931),
            .I(N__40907));
    Span4Mux_h I__8205 (
            .O(N__40928),
            .I(N__40907));
    Span4Mux_h I__8204 (
            .O(N__40925),
            .I(N__40902));
    LocalMux I__8203 (
            .O(N__40922),
            .I(N__40902));
    Span4Mux_v I__8202 (
            .O(N__40919),
            .I(N__40899));
    LocalMux I__8201 (
            .O(N__40916),
            .I(N__40896));
    CEMux I__8200 (
            .O(N__40915),
            .I(N__40893));
    Span4Mux_v I__8199 (
            .O(N__40912),
            .I(N__40888));
    Span4Mux_h I__8198 (
            .O(N__40907),
            .I(N__40888));
    Span4Mux_h I__8197 (
            .O(N__40902),
            .I(N__40885));
    Span4Mux_h I__8196 (
            .O(N__40899),
            .I(N__40878));
    Span4Mux_h I__8195 (
            .O(N__40896),
            .I(N__40878));
    LocalMux I__8194 (
            .O(N__40893),
            .I(N__40878));
    Span4Mux_v I__8193 (
            .O(N__40888),
            .I(N__40875));
    Span4Mux_v I__8192 (
            .O(N__40885),
            .I(N__40872));
    Sp12to4 I__8191 (
            .O(N__40878),
            .I(N__40869));
    Odrv4 I__8190 (
            .O(N__40875),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv4 I__8189 (
            .O(N__40872),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv12 I__8188 (
            .O(N__40869),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    CascadeMux I__8187 (
            .O(N__40862),
            .I(N__40858));
    InMux I__8186 (
            .O(N__40861),
            .I(N__40855));
    InMux I__8185 (
            .O(N__40858),
            .I(N__40852));
    LocalMux I__8184 (
            .O(N__40855),
            .I(N__40846));
    LocalMux I__8183 (
            .O(N__40852),
            .I(N__40846));
    InMux I__8182 (
            .O(N__40851),
            .I(N__40842));
    Span4Mux_v I__8181 (
            .O(N__40846),
            .I(N__40839));
    InMux I__8180 (
            .O(N__40845),
            .I(N__40836));
    LocalMux I__8179 (
            .O(N__40842),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__8178 (
            .O(N__40839),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__8177 (
            .O(N__40836),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__8176 (
            .O(N__40829),
            .I(N__40826));
    LocalMux I__8175 (
            .O(N__40826),
            .I(N__40823));
    Span4Mux_h I__8174 (
            .O(N__40823),
            .I(N__40820));
    Odrv4 I__8173 (
            .O(N__40820),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__8172 (
            .O(N__40817),
            .I(N__40814));
    LocalMux I__8171 (
            .O(N__40814),
            .I(N__40811));
    Span4Mux_h I__8170 (
            .O(N__40811),
            .I(N__40808));
    Odrv4 I__8169 (
            .O(N__40808),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__8168 (
            .O(N__40805),
            .I(N__40801));
    CascadeMux I__8167 (
            .O(N__40804),
            .I(N__40798));
    LocalMux I__8166 (
            .O(N__40801),
            .I(N__40794));
    InMux I__8165 (
            .O(N__40798),
            .I(N__40791));
    InMux I__8164 (
            .O(N__40797),
            .I(N__40788));
    Span4Mux_v I__8163 (
            .O(N__40794),
            .I(N__40783));
    LocalMux I__8162 (
            .O(N__40791),
            .I(N__40783));
    LocalMux I__8161 (
            .O(N__40788),
            .I(N__40780));
    Span4Mux_v I__8160 (
            .O(N__40783),
            .I(N__40776));
    Span4Mux_v I__8159 (
            .O(N__40780),
            .I(N__40773));
    InMux I__8158 (
            .O(N__40779),
            .I(N__40770));
    Odrv4 I__8157 (
            .O(N__40776),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__8156 (
            .O(N__40773),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__8155 (
            .O(N__40770),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__8154 (
            .O(N__40763),
            .I(N__40760));
    LocalMux I__8153 (
            .O(N__40760),
            .I(N__40757));
    Span4Mux_v I__8152 (
            .O(N__40757),
            .I(N__40754));
    Odrv4 I__8151 (
            .O(N__40754),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__8150 (
            .O(N__40751),
            .I(N__40748));
    LocalMux I__8149 (
            .O(N__40748),
            .I(N__40745));
    Span4Mux_h I__8148 (
            .O(N__40745),
            .I(N__40742));
    Odrv4 I__8147 (
            .O(N__40742),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    CascadeMux I__8146 (
            .O(N__40739),
            .I(N__40736));
    InMux I__8145 (
            .O(N__40736),
            .I(N__40729));
    InMux I__8144 (
            .O(N__40735),
            .I(N__40729));
    InMux I__8143 (
            .O(N__40734),
            .I(N__40726));
    LocalMux I__8142 (
            .O(N__40729),
            .I(N__40721));
    LocalMux I__8141 (
            .O(N__40726),
            .I(N__40721));
    Span4Mux_v I__8140 (
            .O(N__40721),
            .I(N__40717));
    InMux I__8139 (
            .O(N__40720),
            .I(N__40714));
    Odrv4 I__8138 (
            .O(N__40717),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__8137 (
            .O(N__40714),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__8136 (
            .O(N__40709),
            .I(N__40706));
    LocalMux I__8135 (
            .O(N__40706),
            .I(N__40703));
    Span4Mux_h I__8134 (
            .O(N__40703),
            .I(N__40700));
    Odrv4 I__8133 (
            .O(N__40700),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__8132 (
            .O(N__40697),
            .I(N__40694));
    LocalMux I__8131 (
            .O(N__40694),
            .I(N__40691));
    Span4Mux_v I__8130 (
            .O(N__40691),
            .I(N__40688));
    Odrv4 I__8129 (
            .O(N__40688),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__8128 (
            .O(N__40685),
            .I(N__40682));
    LocalMux I__8127 (
            .O(N__40682),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    InMux I__8126 (
            .O(N__40679),
            .I(N__40676));
    LocalMux I__8125 (
            .O(N__40676),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ));
    CascadeMux I__8124 (
            .O(N__40673),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ));
    InMux I__8123 (
            .O(N__40670),
            .I(N__40667));
    LocalMux I__8122 (
            .O(N__40667),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    InMux I__8121 (
            .O(N__40664),
            .I(N__40661));
    LocalMux I__8120 (
            .O(N__40661),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    CascadeMux I__8119 (
            .O(N__40658),
            .I(N__40655));
    InMux I__8118 (
            .O(N__40655),
            .I(N__40652));
    LocalMux I__8117 (
            .O(N__40652),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    InMux I__8116 (
            .O(N__40649),
            .I(N__40646));
    LocalMux I__8115 (
            .O(N__40646),
            .I(N__40642));
    InMux I__8114 (
            .O(N__40645),
            .I(N__40639));
    Span4Mux_h I__8113 (
            .O(N__40642),
            .I(N__40636));
    LocalMux I__8112 (
            .O(N__40639),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    Odrv4 I__8111 (
            .O(N__40636),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    InMux I__8110 (
            .O(N__40631),
            .I(N__40611));
    InMux I__8109 (
            .O(N__40630),
            .I(N__40611));
    InMux I__8108 (
            .O(N__40629),
            .I(N__40599));
    InMux I__8107 (
            .O(N__40628),
            .I(N__40599));
    InMux I__8106 (
            .O(N__40627),
            .I(N__40594));
    InMux I__8105 (
            .O(N__40626),
            .I(N__40594));
    InMux I__8104 (
            .O(N__40625),
            .I(N__40589));
    InMux I__8103 (
            .O(N__40624),
            .I(N__40589));
    InMux I__8102 (
            .O(N__40623),
            .I(N__40584));
    InMux I__8101 (
            .O(N__40622),
            .I(N__40584));
    InMux I__8100 (
            .O(N__40621),
            .I(N__40568));
    InMux I__8099 (
            .O(N__40620),
            .I(N__40568));
    InMux I__8098 (
            .O(N__40619),
            .I(N__40568));
    InMux I__8097 (
            .O(N__40618),
            .I(N__40568));
    InMux I__8096 (
            .O(N__40617),
            .I(N__40563));
    InMux I__8095 (
            .O(N__40616),
            .I(N__40563));
    LocalMux I__8094 (
            .O(N__40611),
            .I(N__40560));
    InMux I__8093 (
            .O(N__40610),
            .I(N__40549));
    InMux I__8092 (
            .O(N__40609),
            .I(N__40549));
    InMux I__8091 (
            .O(N__40608),
            .I(N__40549));
    InMux I__8090 (
            .O(N__40607),
            .I(N__40549));
    InMux I__8089 (
            .O(N__40606),
            .I(N__40549));
    InMux I__8088 (
            .O(N__40605),
            .I(N__40544));
    InMux I__8087 (
            .O(N__40604),
            .I(N__40544));
    LocalMux I__8086 (
            .O(N__40599),
            .I(N__40535));
    LocalMux I__8085 (
            .O(N__40594),
            .I(N__40535));
    LocalMux I__8084 (
            .O(N__40589),
            .I(N__40535));
    LocalMux I__8083 (
            .O(N__40584),
            .I(N__40535));
    InMux I__8082 (
            .O(N__40583),
            .I(N__40526));
    InMux I__8081 (
            .O(N__40582),
            .I(N__40526));
    InMux I__8080 (
            .O(N__40581),
            .I(N__40526));
    InMux I__8079 (
            .O(N__40580),
            .I(N__40526));
    InMux I__8078 (
            .O(N__40579),
            .I(N__40519));
    InMux I__8077 (
            .O(N__40578),
            .I(N__40519));
    InMux I__8076 (
            .O(N__40577),
            .I(N__40519));
    LocalMux I__8075 (
            .O(N__40568),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8074 (
            .O(N__40563),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__8073 (
            .O(N__40560),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8072 (
            .O(N__40549),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8071 (
            .O(N__40544),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__8070 (
            .O(N__40535),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8069 (
            .O(N__40526),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__8068 (
            .O(N__40519),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__8067 (
            .O(N__40502),
            .I(N__40499));
    LocalMux I__8066 (
            .O(N__40499),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    CascadeMux I__8065 (
            .O(N__40496),
            .I(elapsed_time_ns_1_RNI35CN9_0_16_cascade_));
    InMux I__8064 (
            .O(N__40493),
            .I(N__40490));
    LocalMux I__8063 (
            .O(N__40490),
            .I(N__40487));
    Span4Mux_h I__8062 (
            .O(N__40487),
            .I(N__40484));
    Odrv4 I__8061 (
            .O(N__40484),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ));
    InMux I__8060 (
            .O(N__40481),
            .I(N__40478));
    LocalMux I__8059 (
            .O(N__40478),
            .I(N__40475));
    Sp12to4 I__8058 (
            .O(N__40475),
            .I(N__40471));
    InMux I__8057 (
            .O(N__40474),
            .I(N__40468));
    Span12Mux_s9_h I__8056 (
            .O(N__40471),
            .I(N__40465));
    LocalMux I__8055 (
            .O(N__40468),
            .I(N__40462));
    Span12Mux_v I__8054 (
            .O(N__40465),
            .I(N__40459));
    Odrv4 I__8053 (
            .O(N__40462),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv12 I__8052 (
            .O(N__40459),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__8051 (
            .O(N__40454),
            .I(N__40451));
    LocalMux I__8050 (
            .O(N__40451),
            .I(N__40447));
    InMux I__8049 (
            .O(N__40450),
            .I(N__40444));
    Span12Mux_s10_h I__8048 (
            .O(N__40447),
            .I(N__40441));
    LocalMux I__8047 (
            .O(N__40444),
            .I(N__40438));
    Span12Mux_v I__8046 (
            .O(N__40441),
            .I(N__40435));
    Odrv4 I__8045 (
            .O(N__40438),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    Odrv12 I__8044 (
            .O(N__40435),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__8043 (
            .O(N__40430),
            .I(N__40427));
    LocalMux I__8042 (
            .O(N__40427),
            .I(N__40424));
    Odrv4 I__8041 (
            .O(N__40424),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_31 ));
    InMux I__8040 (
            .O(N__40421),
            .I(N__40418));
    LocalMux I__8039 (
            .O(N__40418),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ));
    InMux I__8038 (
            .O(N__40415),
            .I(N__40412));
    LocalMux I__8037 (
            .O(N__40412),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    InMux I__8036 (
            .O(N__40409),
            .I(N__40406));
    LocalMux I__8035 (
            .O(N__40406),
            .I(N__40403));
    Span4Mux_h I__8034 (
            .O(N__40403),
            .I(N__40399));
    InMux I__8033 (
            .O(N__40402),
            .I(N__40396));
    Odrv4 I__8032 (
            .O(N__40399),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__8031 (
            .O(N__40396),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__8030 (
            .O(N__40391),
            .I(N__40388));
    LocalMux I__8029 (
            .O(N__40388),
            .I(N__40384));
    CascadeMux I__8028 (
            .O(N__40387),
            .I(N__40381));
    Span4Mux_h I__8027 (
            .O(N__40384),
            .I(N__40378));
    InMux I__8026 (
            .O(N__40381),
            .I(N__40375));
    Odrv4 I__8025 (
            .O(N__40378),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__8024 (
            .O(N__40375),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__8023 (
            .O(N__40370),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ));
    InMux I__8022 (
            .O(N__40367),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ));
    InMux I__8021 (
            .O(N__40364),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ));
    InMux I__8020 (
            .O(N__40361),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ));
    InMux I__8019 (
            .O(N__40358),
            .I(N__40355));
    LocalMux I__8018 (
            .O(N__40355),
            .I(N__40352));
    Span12Mux_s5_h I__8017 (
            .O(N__40352),
            .I(N__40348));
    InMux I__8016 (
            .O(N__40351),
            .I(N__40345));
    Span12Mux_v I__8015 (
            .O(N__40348),
            .I(N__40342));
    LocalMux I__8014 (
            .O(N__40345),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    Odrv12 I__8013 (
            .O(N__40342),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    InMux I__8012 (
            .O(N__40337),
            .I(N__40334));
    LocalMux I__8011 (
            .O(N__40334),
            .I(N__40331));
    Span4Mux_v I__8010 (
            .O(N__40331),
            .I(N__40328));
    Sp12to4 I__8009 (
            .O(N__40328),
            .I(N__40324));
    InMux I__8008 (
            .O(N__40327),
            .I(N__40321));
    Span12Mux_s3_h I__8007 (
            .O(N__40324),
            .I(N__40318));
    LocalMux I__8006 (
            .O(N__40321),
            .I(N__40313));
    Span12Mux_h I__8005 (
            .O(N__40318),
            .I(N__40313));
    Odrv12 I__8004 (
            .O(N__40313),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    InMux I__8003 (
            .O(N__40310),
            .I(N__40307));
    LocalMux I__8002 (
            .O(N__40307),
            .I(N__40304));
    Span4Mux_s3_h I__8001 (
            .O(N__40304),
            .I(N__40301));
    Span4Mux_v I__8000 (
            .O(N__40301),
            .I(N__40297));
    InMux I__7999 (
            .O(N__40300),
            .I(N__40294));
    Sp12to4 I__7998 (
            .O(N__40297),
            .I(N__40291));
    LocalMux I__7997 (
            .O(N__40294),
            .I(N__40286));
    Span12Mux_h I__7996 (
            .O(N__40291),
            .I(N__40286));
    Odrv12 I__7995 (
            .O(N__40286),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__7994 (
            .O(N__40283),
            .I(N__40280));
    LocalMux I__7993 (
            .O(N__40280),
            .I(N__40277));
    Sp12to4 I__7992 (
            .O(N__40277),
            .I(N__40274));
    Span12Mux_s6_h I__7991 (
            .O(N__40274),
            .I(N__40270));
    InMux I__7990 (
            .O(N__40273),
            .I(N__40267));
    Span12Mux_v I__7989 (
            .O(N__40270),
            .I(N__40264));
    LocalMux I__7988 (
            .O(N__40267),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    Odrv12 I__7987 (
            .O(N__40264),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    InMux I__7986 (
            .O(N__40259),
            .I(N__40256));
    LocalMux I__7985 (
            .O(N__40256),
            .I(N__40252));
    InMux I__7984 (
            .O(N__40255),
            .I(N__40249));
    Span12Mux_s8_h I__7983 (
            .O(N__40252),
            .I(N__40246));
    LocalMux I__7982 (
            .O(N__40249),
            .I(N__40243));
    Span12Mux_v I__7981 (
            .O(N__40246),
            .I(N__40240));
    Odrv4 I__7980 (
            .O(N__40243),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    Odrv12 I__7979 (
            .O(N__40240),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    InMux I__7978 (
            .O(N__40235),
            .I(N__40232));
    LocalMux I__7977 (
            .O(N__40232),
            .I(N__40229));
    Span4Mux_h I__7976 (
            .O(N__40229),
            .I(N__40226));
    Span4Mux_h I__7975 (
            .O(N__40226),
            .I(N__40222));
    InMux I__7974 (
            .O(N__40225),
            .I(N__40219));
    Sp12to4 I__7973 (
            .O(N__40222),
            .I(N__40216));
    LocalMux I__7972 (
            .O(N__40219),
            .I(N__40211));
    Span12Mux_v I__7971 (
            .O(N__40216),
            .I(N__40211));
    Odrv12 I__7970 (
            .O(N__40211),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    InMux I__7969 (
            .O(N__40208),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__7968 (
            .O(N__40205),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__7967 (
            .O(N__40202),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__7966 (
            .O(N__40199),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    InMux I__7965 (
            .O(N__40196),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__7964 (
            .O(N__40193),
            .I(bfn_15_24_0_));
    InMux I__7963 (
            .O(N__40190),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__7962 (
            .O(N__40187),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__7961 (
            .O(N__40184),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ));
    InMux I__7960 (
            .O(N__40181),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__7959 (
            .O(N__40178),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__7958 (
            .O(N__40175),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__7957 (
            .O(N__40172),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__7956 (
            .O(N__40169),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__7955 (
            .O(N__40166),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__7954 (
            .O(N__40163),
            .I(bfn_15_23_0_));
    InMux I__7953 (
            .O(N__40160),
            .I(N__40157));
    LocalMux I__7952 (
            .O(N__40157),
            .I(N__40153));
    InMux I__7951 (
            .O(N__40156),
            .I(N__40150));
    Span12Mux_s3_h I__7950 (
            .O(N__40153),
            .I(N__40147));
    LocalMux I__7949 (
            .O(N__40150),
            .I(N__40144));
    Span12Mux_h I__7948 (
            .O(N__40147),
            .I(N__40141));
    Odrv4 I__7947 (
            .O(N__40144),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    Odrv12 I__7946 (
            .O(N__40141),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__7945 (
            .O(N__40136),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__7944 (
            .O(N__40133),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__7943 (
            .O(N__40130),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__7942 (
            .O(N__40127),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__7941 (
            .O(N__40124),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__7940 (
            .O(N__40121),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__7939 (
            .O(N__40118),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__7938 (
            .O(N__40115),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__7937 (
            .O(N__40112),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__7936 (
            .O(N__40109),
            .I(bfn_15_22_0_));
    InMux I__7935 (
            .O(N__40106),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__7934 (
            .O(N__40103),
            .I(N__40100));
    LocalMux I__7933 (
            .O(N__40100),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__7932 (
            .O(N__40097),
            .I(N__40094));
    InMux I__7931 (
            .O(N__40094),
            .I(N__40091));
    LocalMux I__7930 (
            .O(N__40091),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__7929 (
            .O(N__40088),
            .I(N__40085));
    LocalMux I__7928 (
            .O(N__40085),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__7927 (
            .O(N__40082),
            .I(N__40079));
    InMux I__7926 (
            .O(N__40079),
            .I(N__40076));
    LocalMux I__7925 (
            .O(N__40076),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__7924 (
            .O(N__40073),
            .I(N__40070));
    LocalMux I__7923 (
            .O(N__40070),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__7922 (
            .O(N__40067),
            .I(N__40064));
    InMux I__7921 (
            .O(N__40064),
            .I(N__40061));
    LocalMux I__7920 (
            .O(N__40061),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__7919 (
            .O(N__40058),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__7918 (
            .O(N__40055),
            .I(N__40052));
    LocalMux I__7917 (
            .O(N__40052),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    CascadeMux I__7916 (
            .O(N__40049),
            .I(N__40046));
    InMux I__7915 (
            .O(N__40046),
            .I(N__40043));
    LocalMux I__7914 (
            .O(N__40043),
            .I(N__40040));
    Odrv4 I__7913 (
            .O(N__40040),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__7912 (
            .O(N__40037),
            .I(N__40034));
    LocalMux I__7911 (
            .O(N__40034),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__7910 (
            .O(N__40031),
            .I(N__40028));
    InMux I__7909 (
            .O(N__40028),
            .I(N__40025));
    LocalMux I__7908 (
            .O(N__40025),
            .I(N__40022));
    Span4Mux_h I__7907 (
            .O(N__40022),
            .I(N__40019));
    Span4Mux_v I__7906 (
            .O(N__40019),
            .I(N__40016));
    Odrv4 I__7905 (
            .O(N__40016),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__7904 (
            .O(N__40013),
            .I(N__40010));
    LocalMux I__7903 (
            .O(N__40010),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    CascadeMux I__7902 (
            .O(N__40007),
            .I(N__40004));
    InMux I__7901 (
            .O(N__40004),
            .I(N__40001));
    LocalMux I__7900 (
            .O(N__40001),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__7899 (
            .O(N__39998),
            .I(N__39995));
    LocalMux I__7898 (
            .O(N__39995),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__7897 (
            .O(N__39992),
            .I(N__39989));
    InMux I__7896 (
            .O(N__39989),
            .I(N__39986));
    LocalMux I__7895 (
            .O(N__39986),
            .I(N__39983));
    Span4Mux_v I__7894 (
            .O(N__39983),
            .I(N__39980));
    Odrv4 I__7893 (
            .O(N__39980),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__7892 (
            .O(N__39977),
            .I(N__39974));
    LocalMux I__7891 (
            .O(N__39974),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__7890 (
            .O(N__39971),
            .I(N__39968));
    InMux I__7889 (
            .O(N__39968),
            .I(N__39965));
    LocalMux I__7888 (
            .O(N__39965),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    CascadeMux I__7887 (
            .O(N__39962),
            .I(N__39959));
    InMux I__7886 (
            .O(N__39959),
            .I(N__39956));
    LocalMux I__7885 (
            .O(N__39956),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__7884 (
            .O(N__39953),
            .I(N__39950));
    LocalMux I__7883 (
            .O(N__39950),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__7882 (
            .O(N__39947),
            .I(N__39944));
    InMux I__7881 (
            .O(N__39944),
            .I(N__39941));
    LocalMux I__7880 (
            .O(N__39941),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__7879 (
            .O(N__39938),
            .I(N__39935));
    LocalMux I__7878 (
            .O(N__39935),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    CascadeMux I__7877 (
            .O(N__39932),
            .I(N__39929));
    InMux I__7876 (
            .O(N__39929),
            .I(N__39926));
    LocalMux I__7875 (
            .O(N__39926),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__7874 (
            .O(N__39923),
            .I(N__39920));
    LocalMux I__7873 (
            .O(N__39920),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__7872 (
            .O(N__39917),
            .I(N__39914));
    InMux I__7871 (
            .O(N__39914),
            .I(N__39911));
    LocalMux I__7870 (
            .O(N__39911),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__7869 (
            .O(N__39908),
            .I(N__39905));
    LocalMux I__7868 (
            .O(N__39905),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    InMux I__7867 (
            .O(N__39902),
            .I(N__39898));
    InMux I__7866 (
            .O(N__39901),
            .I(N__39894));
    LocalMux I__7865 (
            .O(N__39898),
            .I(N__39891));
    InMux I__7864 (
            .O(N__39897),
            .I(N__39888));
    LocalMux I__7863 (
            .O(N__39894),
            .I(N__39885));
    Span4Mux_v I__7862 (
            .O(N__39891),
            .I(N__39882));
    LocalMux I__7861 (
            .O(N__39888),
            .I(N__39877));
    Span4Mux_v I__7860 (
            .O(N__39885),
            .I(N__39877));
    Odrv4 I__7859 (
            .O(N__39882),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__7858 (
            .O(N__39877),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__7857 (
            .O(N__39872),
            .I(N__39868));
    InMux I__7856 (
            .O(N__39871),
            .I(N__39865));
    LocalMux I__7855 (
            .O(N__39868),
            .I(N__39862));
    LocalMux I__7854 (
            .O(N__39865),
            .I(N__39859));
    Span4Mux_h I__7853 (
            .O(N__39862),
            .I(N__39856));
    Span4Mux_h I__7852 (
            .O(N__39859),
            .I(N__39853));
    Odrv4 I__7851 (
            .O(N__39856),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv4 I__7850 (
            .O(N__39853),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    CascadeMux I__7849 (
            .O(N__39848),
            .I(N__39845));
    InMux I__7848 (
            .O(N__39845),
            .I(N__39842));
    LocalMux I__7847 (
            .O(N__39842),
            .I(N__39839));
    Odrv4 I__7846 (
            .O(N__39839),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__7845 (
            .O(N__39836),
            .I(N__39833));
    LocalMux I__7844 (
            .O(N__39833),
            .I(N__39830));
    Odrv4 I__7843 (
            .O(N__39830),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__7842 (
            .O(N__39827),
            .I(N__39824));
    InMux I__7841 (
            .O(N__39824),
            .I(N__39821));
    LocalMux I__7840 (
            .O(N__39821),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__7839 (
            .O(N__39818),
            .I(N__39815));
    LocalMux I__7838 (
            .O(N__39815),
            .I(N__39812));
    Odrv12 I__7837 (
            .O(N__39812),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__7836 (
            .O(N__39809),
            .I(N__39806));
    InMux I__7835 (
            .O(N__39806),
            .I(N__39803));
    LocalMux I__7834 (
            .O(N__39803),
            .I(N__39800));
    Odrv4 I__7833 (
            .O(N__39800),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__7832 (
            .O(N__39797),
            .I(N__39794));
    LocalMux I__7831 (
            .O(N__39794),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__7830 (
            .O(N__39791),
            .I(N__39788));
    InMux I__7829 (
            .O(N__39788),
            .I(N__39785));
    LocalMux I__7828 (
            .O(N__39785),
            .I(N__39782));
    Odrv12 I__7827 (
            .O(N__39782),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__7826 (
            .O(N__39779),
            .I(N__39774));
    InMux I__7825 (
            .O(N__39778),
            .I(N__39771));
    InMux I__7824 (
            .O(N__39777),
            .I(N__39768));
    InMux I__7823 (
            .O(N__39774),
            .I(N__39765));
    LocalMux I__7822 (
            .O(N__39771),
            .I(N__39762));
    LocalMux I__7821 (
            .O(N__39768),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__7820 (
            .O(N__39765),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__7819 (
            .O(N__39762),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__7818 (
            .O(N__39755),
            .I(N__39750));
    InMux I__7817 (
            .O(N__39754),
            .I(N__39747));
    InMux I__7816 (
            .O(N__39753),
            .I(N__39744));
    LocalMux I__7815 (
            .O(N__39750),
            .I(N__39739));
    LocalMux I__7814 (
            .O(N__39747),
            .I(N__39739));
    LocalMux I__7813 (
            .O(N__39744),
            .I(N__39733));
    Span4Mux_v I__7812 (
            .O(N__39739),
            .I(N__39733));
    InMux I__7811 (
            .O(N__39738),
            .I(N__39730));
    Odrv4 I__7810 (
            .O(N__39733),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__7809 (
            .O(N__39730),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    CascadeMux I__7808 (
            .O(N__39725),
            .I(N__39721));
    CascadeMux I__7807 (
            .O(N__39724),
            .I(N__39718));
    InMux I__7806 (
            .O(N__39721),
            .I(N__39715));
    InMux I__7805 (
            .O(N__39718),
            .I(N__39712));
    LocalMux I__7804 (
            .O(N__39715),
            .I(N__39709));
    LocalMux I__7803 (
            .O(N__39712),
            .I(N__39703));
    Span4Mux_h I__7802 (
            .O(N__39709),
            .I(N__39703));
    InMux I__7801 (
            .O(N__39708),
            .I(N__39700));
    Span4Mux_v I__7800 (
            .O(N__39703),
            .I(N__39696));
    LocalMux I__7799 (
            .O(N__39700),
            .I(N__39693));
    InMux I__7798 (
            .O(N__39699),
            .I(N__39690));
    Odrv4 I__7797 (
            .O(N__39696),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv12 I__7796 (
            .O(N__39693),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__7795 (
            .O(N__39690),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__7794 (
            .O(N__39683),
            .I(N__39678));
    InMux I__7793 (
            .O(N__39682),
            .I(N__39675));
    InMux I__7792 (
            .O(N__39681),
            .I(N__39672));
    LocalMux I__7791 (
            .O(N__39678),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__7790 (
            .O(N__39675),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__7789 (
            .O(N__39672),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__7788 (
            .O(N__39665),
            .I(N__39661));
    InMux I__7787 (
            .O(N__39664),
            .I(N__39643));
    InMux I__7786 (
            .O(N__39661),
            .I(N__39643));
    InMux I__7785 (
            .O(N__39660),
            .I(N__39640));
    InMux I__7784 (
            .O(N__39659),
            .I(N__39628));
    InMux I__7783 (
            .O(N__39658),
            .I(N__39628));
    InMux I__7782 (
            .O(N__39657),
            .I(N__39615));
    InMux I__7781 (
            .O(N__39656),
            .I(N__39615));
    InMux I__7780 (
            .O(N__39655),
            .I(N__39615));
    InMux I__7779 (
            .O(N__39654),
            .I(N__39615));
    InMux I__7778 (
            .O(N__39653),
            .I(N__39615));
    InMux I__7777 (
            .O(N__39652),
            .I(N__39615));
    InMux I__7776 (
            .O(N__39651),
            .I(N__39606));
    InMux I__7775 (
            .O(N__39650),
            .I(N__39606));
    InMux I__7774 (
            .O(N__39649),
            .I(N__39606));
    InMux I__7773 (
            .O(N__39648),
            .I(N__39606));
    LocalMux I__7772 (
            .O(N__39643),
            .I(N__39601));
    LocalMux I__7771 (
            .O(N__39640),
            .I(N__39601));
    InMux I__7770 (
            .O(N__39639),
            .I(N__39586));
    InMux I__7769 (
            .O(N__39638),
            .I(N__39586));
    InMux I__7768 (
            .O(N__39637),
            .I(N__39586));
    InMux I__7767 (
            .O(N__39636),
            .I(N__39586));
    InMux I__7766 (
            .O(N__39635),
            .I(N__39586));
    InMux I__7765 (
            .O(N__39634),
            .I(N__39586));
    InMux I__7764 (
            .O(N__39633),
            .I(N__39586));
    LocalMux I__7763 (
            .O(N__39628),
            .I(N__39582));
    LocalMux I__7762 (
            .O(N__39615),
            .I(N__39579));
    LocalMux I__7761 (
            .O(N__39606),
            .I(N__39574));
    Span4Mux_v I__7760 (
            .O(N__39601),
            .I(N__39569));
    LocalMux I__7759 (
            .O(N__39586),
            .I(N__39569));
    InMux I__7758 (
            .O(N__39585),
            .I(N__39566));
    Span4Mux_v I__7757 (
            .O(N__39582),
            .I(N__39563));
    Span4Mux_h I__7756 (
            .O(N__39579),
            .I(N__39560));
    InMux I__7755 (
            .O(N__39578),
            .I(N__39555));
    InMux I__7754 (
            .O(N__39577),
            .I(N__39555));
    Span4Mux_h I__7753 (
            .O(N__39574),
            .I(N__39552));
    Odrv4 I__7752 (
            .O(N__39569),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__7751 (
            .O(N__39566),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__7750 (
            .O(N__39563),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__7749 (
            .O(N__39560),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__7748 (
            .O(N__39555),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__7747 (
            .O(N__39552),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__7746 (
            .O(N__39539),
            .I(N__39534));
    InMux I__7745 (
            .O(N__39538),
            .I(N__39531));
    InMux I__7744 (
            .O(N__39537),
            .I(N__39528));
    InMux I__7743 (
            .O(N__39534),
            .I(N__39525));
    LocalMux I__7742 (
            .O(N__39531),
            .I(N__39522));
    LocalMux I__7741 (
            .O(N__39528),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__7740 (
            .O(N__39525),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__7739 (
            .O(N__39522),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__7738 (
            .O(N__39515),
            .I(N__39510));
    InMux I__7737 (
            .O(N__39514),
            .I(N__39507));
    InMux I__7736 (
            .O(N__39513),
            .I(N__39504));
    LocalMux I__7735 (
            .O(N__39510),
            .I(N__39501));
    LocalMux I__7734 (
            .O(N__39507),
            .I(N__39496));
    LocalMux I__7733 (
            .O(N__39504),
            .I(N__39496));
    Span4Mux_v I__7732 (
            .O(N__39501),
            .I(N__39490));
    Span4Mux_v I__7731 (
            .O(N__39496),
            .I(N__39490));
    InMux I__7730 (
            .O(N__39495),
            .I(N__39487));
    Odrv4 I__7729 (
            .O(N__39490),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__7728 (
            .O(N__39487),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    CascadeMux I__7727 (
            .O(N__39482),
            .I(N__39477));
    InMux I__7726 (
            .O(N__39481),
            .I(N__39474));
    InMux I__7725 (
            .O(N__39480),
            .I(N__39471));
    InMux I__7724 (
            .O(N__39477),
            .I(N__39468));
    LocalMux I__7723 (
            .O(N__39474),
            .I(N__39463));
    LocalMux I__7722 (
            .O(N__39471),
            .I(N__39463));
    LocalMux I__7721 (
            .O(N__39468),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__7720 (
            .O(N__39463),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__7719 (
            .O(N__39458),
            .I(N__39455));
    LocalMux I__7718 (
            .O(N__39455),
            .I(N__39452));
    Span4Mux_v I__7717 (
            .O(N__39452),
            .I(N__39447));
    InMux I__7716 (
            .O(N__39451),
            .I(N__39444));
    InMux I__7715 (
            .O(N__39450),
            .I(N__39441));
    Span4Mux_h I__7714 (
            .O(N__39447),
            .I(N__39436));
    LocalMux I__7713 (
            .O(N__39444),
            .I(N__39436));
    LocalMux I__7712 (
            .O(N__39441),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__7711 (
            .O(N__39436),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__7710 (
            .O(N__39431),
            .I(N__39426));
    InMux I__7709 (
            .O(N__39430),
            .I(N__39423));
    CascadeMux I__7708 (
            .O(N__39429),
            .I(N__39420));
    LocalMux I__7707 (
            .O(N__39426),
            .I(N__39414));
    LocalMux I__7706 (
            .O(N__39423),
            .I(N__39414));
    InMux I__7705 (
            .O(N__39420),
            .I(N__39411));
    InMux I__7704 (
            .O(N__39419),
            .I(N__39408));
    Span4Mux_v I__7703 (
            .O(N__39414),
            .I(N__39405));
    LocalMux I__7702 (
            .O(N__39411),
            .I(N__39400));
    LocalMux I__7701 (
            .O(N__39408),
            .I(N__39400));
    Span4Mux_v I__7700 (
            .O(N__39405),
            .I(N__39397));
    Span4Mux_h I__7699 (
            .O(N__39400),
            .I(N__39394));
    Odrv4 I__7698 (
            .O(N__39397),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__7697 (
            .O(N__39394),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    CascadeMux I__7696 (
            .O(N__39389),
            .I(N__39386));
    InMux I__7695 (
            .O(N__39386),
            .I(N__39382));
    InMux I__7694 (
            .O(N__39385),
            .I(N__39378));
    LocalMux I__7693 (
            .O(N__39382),
            .I(N__39375));
    InMux I__7692 (
            .O(N__39381),
            .I(N__39372));
    LocalMux I__7691 (
            .O(N__39378),
            .I(N__39369));
    Span4Mux_h I__7690 (
            .O(N__39375),
            .I(N__39364));
    LocalMux I__7689 (
            .O(N__39372),
            .I(N__39364));
    Span4Mux_v I__7688 (
            .O(N__39369),
            .I(N__39358));
    Span4Mux_v I__7687 (
            .O(N__39364),
            .I(N__39358));
    InMux I__7686 (
            .O(N__39363),
            .I(N__39355));
    Odrv4 I__7685 (
            .O(N__39358),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__7684 (
            .O(N__39355),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__7683 (
            .O(N__39350),
            .I(N__39343));
    InMux I__7682 (
            .O(N__39349),
            .I(N__39343));
    InMux I__7681 (
            .O(N__39348),
            .I(N__39340));
    LocalMux I__7680 (
            .O(N__39343),
            .I(N__39336));
    LocalMux I__7679 (
            .O(N__39340),
            .I(N__39333));
    InMux I__7678 (
            .O(N__39339),
            .I(N__39330));
    Span4Mux_h I__7677 (
            .O(N__39336),
            .I(N__39327));
    Sp12to4 I__7676 (
            .O(N__39333),
            .I(N__39322));
    LocalMux I__7675 (
            .O(N__39330),
            .I(N__39322));
    Odrv4 I__7674 (
            .O(N__39327),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv12 I__7673 (
            .O(N__39322),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__7672 (
            .O(N__39317),
            .I(N__39314));
    LocalMux I__7671 (
            .O(N__39314),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__7670 (
            .O(N__39311),
            .I(N__39308));
    LocalMux I__7669 (
            .O(N__39308),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__7668 (
            .O(N__39305),
            .I(N__39302));
    InMux I__7667 (
            .O(N__39302),
            .I(N__39298));
    InMux I__7666 (
            .O(N__39301),
            .I(N__39294));
    LocalMux I__7665 (
            .O(N__39298),
            .I(N__39291));
    InMux I__7664 (
            .O(N__39297),
            .I(N__39288));
    LocalMux I__7663 (
            .O(N__39294),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__7662 (
            .O(N__39291),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__7661 (
            .O(N__39288),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__7660 (
            .O(N__39281),
            .I(N__39276));
    InMux I__7659 (
            .O(N__39280),
            .I(N__39273));
    InMux I__7658 (
            .O(N__39279),
            .I(N__39270));
    LocalMux I__7657 (
            .O(N__39276),
            .I(N__39267));
    LocalMux I__7656 (
            .O(N__39273),
            .I(N__39264));
    LocalMux I__7655 (
            .O(N__39270),
            .I(N__39260));
    Span4Mux_v I__7654 (
            .O(N__39267),
            .I(N__39257));
    Span4Mux_v I__7653 (
            .O(N__39264),
            .I(N__39254));
    InMux I__7652 (
            .O(N__39263),
            .I(N__39251));
    Odrv12 I__7651 (
            .O(N__39260),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__7650 (
            .O(N__39257),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__7649 (
            .O(N__39254),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__7648 (
            .O(N__39251),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    CascadeMux I__7647 (
            .O(N__39242),
            .I(N__39237));
    InMux I__7646 (
            .O(N__39241),
            .I(N__39234));
    InMux I__7645 (
            .O(N__39240),
            .I(N__39231));
    InMux I__7644 (
            .O(N__39237),
            .I(N__39228));
    LocalMux I__7643 (
            .O(N__39234),
            .I(N__39223));
    LocalMux I__7642 (
            .O(N__39231),
            .I(N__39223));
    LocalMux I__7641 (
            .O(N__39228),
            .I(\current_shift_inst.un4_control_input1_21 ));
    Odrv4 I__7640 (
            .O(N__39223),
            .I(\current_shift_inst.un4_control_input1_21 ));
    CascadeMux I__7639 (
            .O(N__39218),
            .I(N__39215));
    InMux I__7638 (
            .O(N__39215),
            .I(N__39210));
    InMux I__7637 (
            .O(N__39214),
            .I(N__39207));
    InMux I__7636 (
            .O(N__39213),
            .I(N__39204));
    LocalMux I__7635 (
            .O(N__39210),
            .I(N__39201));
    LocalMux I__7634 (
            .O(N__39207),
            .I(N__39198));
    LocalMux I__7633 (
            .O(N__39204),
            .I(N__39191));
    Span4Mux_v I__7632 (
            .O(N__39201),
            .I(N__39191));
    Span4Mux_v I__7631 (
            .O(N__39198),
            .I(N__39191));
    Span4Mux_v I__7630 (
            .O(N__39191),
            .I(N__39187));
    InMux I__7629 (
            .O(N__39190),
            .I(N__39184));
    Odrv4 I__7628 (
            .O(N__39187),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__7627 (
            .O(N__39184),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__7626 (
            .O(N__39179),
            .I(N__39175));
    CascadeMux I__7625 (
            .O(N__39178),
            .I(N__39171));
    LocalMux I__7624 (
            .O(N__39175),
            .I(N__39168));
    InMux I__7623 (
            .O(N__39174),
            .I(N__39165));
    InMux I__7622 (
            .O(N__39171),
            .I(N__39162));
    Span4Mux_v I__7621 (
            .O(N__39168),
            .I(N__39159));
    LocalMux I__7620 (
            .O(N__39165),
            .I(N__39156));
    LocalMux I__7619 (
            .O(N__39162),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__7618 (
            .O(N__39159),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__7617 (
            .O(N__39156),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__7616 (
            .O(N__39149),
            .I(N__39144));
    InMux I__7615 (
            .O(N__39148),
            .I(N__39141));
    InMux I__7614 (
            .O(N__39147),
            .I(N__39138));
    LocalMux I__7613 (
            .O(N__39144),
            .I(N__39135));
    LocalMux I__7612 (
            .O(N__39141),
            .I(N__39130));
    LocalMux I__7611 (
            .O(N__39138),
            .I(N__39130));
    Span4Mux_h I__7610 (
            .O(N__39135),
            .I(N__39124));
    Span4Mux_v I__7609 (
            .O(N__39130),
            .I(N__39124));
    InMux I__7608 (
            .O(N__39129),
            .I(N__39121));
    Odrv4 I__7607 (
            .O(N__39124),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__7606 (
            .O(N__39121),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__7605 (
            .O(N__39116),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__7604 (
            .O(N__39113),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__7603 (
            .O(N__39110),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__7602 (
            .O(N__39107),
            .I(N__39104));
    LocalMux I__7601 (
            .O(N__39104),
            .I(N__39100));
    InMux I__7600 (
            .O(N__39103),
            .I(N__39097));
    Span4Mux_h I__7599 (
            .O(N__39100),
            .I(N__39093));
    LocalMux I__7598 (
            .O(N__39097),
            .I(N__39090));
    InMux I__7597 (
            .O(N__39096),
            .I(N__39087));
    Odrv4 I__7596 (
            .O(N__39093),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__7595 (
            .O(N__39090),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    LocalMux I__7594 (
            .O(N__39087),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CEMux I__7593 (
            .O(N__39080),
            .I(N__39059));
    CEMux I__7592 (
            .O(N__39079),
            .I(N__39059));
    CEMux I__7591 (
            .O(N__39078),
            .I(N__39059));
    CEMux I__7590 (
            .O(N__39077),
            .I(N__39059));
    CEMux I__7589 (
            .O(N__39076),
            .I(N__39059));
    CEMux I__7588 (
            .O(N__39075),
            .I(N__39059));
    CEMux I__7587 (
            .O(N__39074),
            .I(N__39059));
    GlobalMux I__7586 (
            .O(N__39059),
            .I(N__39056));
    gio2CtrlBuf I__7585 (
            .O(N__39056),
            .I(\current_shift_inst.timer_s1.N_163_i_g ));
    CascadeMux I__7584 (
            .O(N__39053),
            .I(N__39050));
    InMux I__7583 (
            .O(N__39050),
            .I(N__39046));
    InMux I__7582 (
            .O(N__39049),
            .I(N__39043));
    LocalMux I__7581 (
            .O(N__39046),
            .I(N__39039));
    LocalMux I__7580 (
            .O(N__39043),
            .I(N__39036));
    InMux I__7579 (
            .O(N__39042),
            .I(N__39033));
    Span4Mux_h I__7578 (
            .O(N__39039),
            .I(N__39029));
    Span4Mux_h I__7577 (
            .O(N__39036),
            .I(N__39026));
    LocalMux I__7576 (
            .O(N__39033),
            .I(N__39023));
    InMux I__7575 (
            .O(N__39032),
            .I(N__39020));
    Odrv4 I__7574 (
            .O(N__39029),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__7573 (
            .O(N__39026),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv12 I__7572 (
            .O(N__39023),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__7571 (
            .O(N__39020),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__7570 (
            .O(N__39011),
            .I(N__39007));
    InMux I__7569 (
            .O(N__39010),
            .I(N__39003));
    LocalMux I__7568 (
            .O(N__39007),
            .I(N__39000));
    InMux I__7567 (
            .O(N__39006),
            .I(N__38997));
    LocalMux I__7566 (
            .O(N__39003),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__7565 (
            .O(N__39000),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__7564 (
            .O(N__38997),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__7563 (
            .O(N__38990),
            .I(N__38983));
    InMux I__7562 (
            .O(N__38989),
            .I(N__38983));
    InMux I__7561 (
            .O(N__38988),
            .I(N__38980));
    LocalMux I__7560 (
            .O(N__38983),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__7559 (
            .O(N__38980),
            .I(\current_shift_inst.un4_control_input1_6 ));
    CascadeMux I__7558 (
            .O(N__38975),
            .I(N__38971));
    InMux I__7557 (
            .O(N__38974),
            .I(N__38966));
    InMux I__7556 (
            .O(N__38971),
            .I(N__38966));
    LocalMux I__7555 (
            .O(N__38966),
            .I(N__38962));
    InMux I__7554 (
            .O(N__38965),
            .I(N__38959));
    Span4Mux_v I__7553 (
            .O(N__38962),
            .I(N__38956));
    LocalMux I__7552 (
            .O(N__38959),
            .I(N__38953));
    Span4Mux_h I__7551 (
            .O(N__38956),
            .I(N__38949));
    Span4Mux_v I__7550 (
            .O(N__38953),
            .I(N__38946));
    InMux I__7549 (
            .O(N__38952),
            .I(N__38943));
    Odrv4 I__7548 (
            .O(N__38949),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__7547 (
            .O(N__38946),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__7546 (
            .O(N__38943),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__7545 (
            .O(N__38936),
            .I(N__38930));
    InMux I__7544 (
            .O(N__38935),
            .I(N__38930));
    LocalMux I__7543 (
            .O(N__38930),
            .I(N__38926));
    InMux I__7542 (
            .O(N__38929),
            .I(N__38923));
    Span4Mux_v I__7541 (
            .O(N__38926),
            .I(N__38919));
    LocalMux I__7540 (
            .O(N__38923),
            .I(N__38916));
    InMux I__7539 (
            .O(N__38922),
            .I(N__38913));
    Odrv4 I__7538 (
            .O(N__38919),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv12 I__7537 (
            .O(N__38916),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__7536 (
            .O(N__38913),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    CascadeMux I__7535 (
            .O(N__38906),
            .I(N__38903));
    InMux I__7534 (
            .O(N__38903),
            .I(N__38896));
    InMux I__7533 (
            .O(N__38902),
            .I(N__38896));
    InMux I__7532 (
            .O(N__38901),
            .I(N__38893));
    LocalMux I__7531 (
            .O(N__38896),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__7530 (
            .O(N__38893),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__7529 (
            .O(N__38888),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__7528 (
            .O(N__38885),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__7527 (
            .O(N__38882),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__7526 (
            .O(N__38879),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__7525 (
            .O(N__38876),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__7524 (
            .O(N__38873),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__7523 (
            .O(N__38870),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__7522 (
            .O(N__38867),
            .I(N__38860));
    InMux I__7521 (
            .O(N__38866),
            .I(N__38860));
    InMux I__7520 (
            .O(N__38865),
            .I(N__38856));
    LocalMux I__7519 (
            .O(N__38860),
            .I(N__38853));
    InMux I__7518 (
            .O(N__38859),
            .I(N__38850));
    LocalMux I__7517 (
            .O(N__38856),
            .I(N__38847));
    Span4Mux_v I__7516 (
            .O(N__38853),
            .I(N__38842));
    LocalMux I__7515 (
            .O(N__38850),
            .I(N__38842));
    Sp12to4 I__7514 (
            .O(N__38847),
            .I(N__38839));
    Span4Mux_v I__7513 (
            .O(N__38842),
            .I(N__38836));
    Odrv12 I__7512 (
            .O(N__38839),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__7511 (
            .O(N__38836),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__7510 (
            .O(N__38831),
            .I(bfn_15_13_0_));
    InMux I__7509 (
            .O(N__38828),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__7508 (
            .O(N__38825),
            .I(bfn_15_11_0_));
    CascadeMux I__7507 (
            .O(N__38822),
            .I(N__38818));
    CascadeMux I__7506 (
            .O(N__38821),
            .I(N__38815));
    InMux I__7505 (
            .O(N__38818),
            .I(N__38812));
    InMux I__7504 (
            .O(N__38815),
            .I(N__38809));
    LocalMux I__7503 (
            .O(N__38812),
            .I(N__38805));
    LocalMux I__7502 (
            .O(N__38809),
            .I(N__38802));
    InMux I__7501 (
            .O(N__38808),
            .I(N__38799));
    Span4Mux_h I__7500 (
            .O(N__38805),
            .I(N__38794));
    Span4Mux_h I__7499 (
            .O(N__38802),
            .I(N__38794));
    LocalMux I__7498 (
            .O(N__38799),
            .I(N__38791));
    Span4Mux_v I__7497 (
            .O(N__38794),
            .I(N__38787));
    Span4Mux_v I__7496 (
            .O(N__38791),
            .I(N__38784));
    InMux I__7495 (
            .O(N__38790),
            .I(N__38781));
    Odrv4 I__7494 (
            .O(N__38787),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__7493 (
            .O(N__38784),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__7492 (
            .O(N__38781),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__7491 (
            .O(N__38774),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__7490 (
            .O(N__38771),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__7489 (
            .O(N__38768),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__7488 (
            .O(N__38765),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__7487 (
            .O(N__38762),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7486 (
            .O(N__38759),
            .I(N__38756));
    InMux I__7485 (
            .O(N__38756),
            .I(N__38753));
    LocalMux I__7484 (
            .O(N__38753),
            .I(N__38748));
    InMux I__7483 (
            .O(N__38752),
            .I(N__38745));
    InMux I__7482 (
            .O(N__38751),
            .I(N__38742));
    Span4Mux_h I__7481 (
            .O(N__38748),
            .I(N__38737));
    LocalMux I__7480 (
            .O(N__38745),
            .I(N__38737));
    LocalMux I__7479 (
            .O(N__38742),
            .I(N__38734));
    Span4Mux_v I__7478 (
            .O(N__38737),
            .I(N__38731));
    Span4Mux_h I__7477 (
            .O(N__38734),
            .I(N__38727));
    Span4Mux_v I__7476 (
            .O(N__38731),
            .I(N__38724));
    InMux I__7475 (
            .O(N__38730),
            .I(N__38721));
    Odrv4 I__7474 (
            .O(N__38727),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__7473 (
            .O(N__38724),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__7472 (
            .O(N__38721),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__7471 (
            .O(N__38714),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__7470 (
            .O(N__38711),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__7469 (
            .O(N__38708),
            .I(bfn_15_12_0_));
    InMux I__7468 (
            .O(N__38705),
            .I(N__38701));
    InMux I__7467 (
            .O(N__38704),
            .I(N__38698));
    LocalMux I__7466 (
            .O(N__38701),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    LocalMux I__7465 (
            .O(N__38698),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__7464 (
            .O(N__38693),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__7463 (
            .O(N__38690),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__7462 (
            .O(N__38687),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__7461 (
            .O(N__38684),
            .I(N__38680));
    InMux I__7460 (
            .O(N__38683),
            .I(N__38677));
    InMux I__7459 (
            .O(N__38680),
            .I(N__38674));
    LocalMux I__7458 (
            .O(N__38677),
            .I(N__38670));
    LocalMux I__7457 (
            .O(N__38674),
            .I(N__38667));
    InMux I__7456 (
            .O(N__38673),
            .I(N__38664));
    Span4Mux_h I__7455 (
            .O(N__38670),
            .I(N__38659));
    Span4Mux_h I__7454 (
            .O(N__38667),
            .I(N__38659));
    LocalMux I__7453 (
            .O(N__38664),
            .I(N__38656));
    Span4Mux_v I__7452 (
            .O(N__38659),
            .I(N__38652));
    Span4Mux_v I__7451 (
            .O(N__38656),
            .I(N__38649));
    InMux I__7450 (
            .O(N__38655),
            .I(N__38646));
    Odrv4 I__7449 (
            .O(N__38652),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__7448 (
            .O(N__38649),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__7447 (
            .O(N__38646),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__7446 (
            .O(N__38639),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__7445 (
            .O(N__38636),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__7444 (
            .O(N__38633),
            .I(N__38630));
    InMux I__7443 (
            .O(N__38630),
            .I(N__38626));
    InMux I__7442 (
            .O(N__38629),
            .I(N__38622));
    LocalMux I__7441 (
            .O(N__38626),
            .I(N__38619));
    InMux I__7440 (
            .O(N__38625),
            .I(N__38616));
    LocalMux I__7439 (
            .O(N__38622),
            .I(N__38613));
    Sp12to4 I__7438 (
            .O(N__38619),
            .I(N__38608));
    LocalMux I__7437 (
            .O(N__38616),
            .I(N__38608));
    Span4Mux_v I__7436 (
            .O(N__38613),
            .I(N__38605));
    Span12Mux_v I__7435 (
            .O(N__38608),
            .I(N__38601));
    Span4Mux_v I__7434 (
            .O(N__38605),
            .I(N__38598));
    InMux I__7433 (
            .O(N__38604),
            .I(N__38595));
    Odrv12 I__7432 (
            .O(N__38601),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__7431 (
            .O(N__38598),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__7430 (
            .O(N__38595),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__7429 (
            .O(N__38588),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__7428 (
            .O(N__38585),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__7427 (
            .O(N__38582),
            .I(N__38578));
    InMux I__7426 (
            .O(N__38581),
            .I(N__38575));
    LocalMux I__7425 (
            .O(N__38578),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__7424 (
            .O(N__38575),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    InMux I__7423 (
            .O(N__38570),
            .I(N__38566));
    InMux I__7422 (
            .O(N__38569),
            .I(N__38563));
    LocalMux I__7421 (
            .O(N__38566),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    LocalMux I__7420 (
            .O(N__38563),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    InMux I__7419 (
            .O(N__38558),
            .I(N__38555));
    LocalMux I__7418 (
            .O(N__38555),
            .I(N__38552));
    Span4Mux_v I__7417 (
            .O(N__38552),
            .I(N__38548));
    InMux I__7416 (
            .O(N__38551),
            .I(N__38545));
    Span4Mux_h I__7415 (
            .O(N__38548),
            .I(N__38542));
    LocalMux I__7414 (
            .O(N__38545),
            .I(N__38539));
    Span4Mux_h I__7413 (
            .O(N__38542),
            .I(N__38534));
    Span4Mux_v I__7412 (
            .O(N__38539),
            .I(N__38534));
    Span4Mux_v I__7411 (
            .O(N__38534),
            .I(N__38529));
    InMux I__7410 (
            .O(N__38533),
            .I(N__38526));
    InMux I__7409 (
            .O(N__38532),
            .I(N__38523));
    Span4Mux_v I__7408 (
            .O(N__38529),
            .I(N__38520));
    LocalMux I__7407 (
            .O(N__38526),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__7406 (
            .O(N__38523),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__7405 (
            .O(N__38520),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__7404 (
            .O(N__38513),
            .I(N__38509));
    InMux I__7403 (
            .O(N__38512),
            .I(N__38506));
    LocalMux I__7402 (
            .O(N__38509),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__7401 (
            .O(N__38506),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__7400 (
            .O(N__38501),
            .I(N__38498));
    LocalMux I__7399 (
            .O(N__38498),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    CascadeMux I__7398 (
            .O(N__38495),
            .I(elapsed_time_ns_1_RNI25DN9_0_24_cascade_));
    InMux I__7397 (
            .O(N__38492),
            .I(N__38489));
    LocalMux I__7396 (
            .O(N__38489),
            .I(N__38486));
    Span4Mux_h I__7395 (
            .O(N__38486),
            .I(N__38483));
    Odrv4 I__7394 (
            .O(N__38483),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ));
    InMux I__7393 (
            .O(N__38480),
            .I(N__38476));
    InMux I__7392 (
            .O(N__38479),
            .I(N__38473));
    LocalMux I__7391 (
            .O(N__38476),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    LocalMux I__7390 (
            .O(N__38473),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    InMux I__7389 (
            .O(N__38468),
            .I(N__38465));
    LocalMux I__7388 (
            .O(N__38465),
            .I(N__38462));
    Span4Mux_h I__7387 (
            .O(N__38462),
            .I(N__38459));
    Odrv4 I__7386 (
            .O(N__38459),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ));
    InMux I__7385 (
            .O(N__38456),
            .I(N__38452));
    InMux I__7384 (
            .O(N__38455),
            .I(N__38449));
    LocalMux I__7383 (
            .O(N__38452),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__7382 (
            .O(N__38449),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    CascadeMux I__7381 (
            .O(N__38444),
            .I(elapsed_time_ns_1_RNIG23T9_0_4_cascade_));
    InMux I__7380 (
            .O(N__38441),
            .I(N__38438));
    LocalMux I__7379 (
            .O(N__38438),
            .I(N__38435));
    Span4Mux_h I__7378 (
            .O(N__38435),
            .I(N__38432));
    Odrv4 I__7377 (
            .O(N__38432),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ));
    InMux I__7376 (
            .O(N__38429),
            .I(N__38426));
    LocalMux I__7375 (
            .O(N__38426),
            .I(N__38422));
    InMux I__7374 (
            .O(N__38425),
            .I(N__38419));
    Span4Mux_v I__7373 (
            .O(N__38422),
            .I(N__38416));
    LocalMux I__7372 (
            .O(N__38419),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv4 I__7371 (
            .O(N__38416),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    CascadeMux I__7370 (
            .O(N__38411),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27_cascade_ ));
    InMux I__7369 (
            .O(N__38408),
            .I(N__38405));
    LocalMux I__7368 (
            .O(N__38405),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    CascadeMux I__7367 (
            .O(N__38402),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    InMux I__7366 (
            .O(N__38399),
            .I(N__38395));
    InMux I__7365 (
            .O(N__38398),
            .I(N__38392));
    LocalMux I__7364 (
            .O(N__38395),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    LocalMux I__7363 (
            .O(N__38392),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__7362 (
            .O(N__38387),
            .I(N__38383));
    InMux I__7361 (
            .O(N__38386),
            .I(N__38380));
    LocalMux I__7360 (
            .O(N__38383),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    LocalMux I__7359 (
            .O(N__38380),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    InMux I__7358 (
            .O(N__38375),
            .I(N__38372));
    LocalMux I__7357 (
            .O(N__38372),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    CascadeMux I__7356 (
            .O(N__38369),
            .I(elapsed_time_ns_1_RNI13CN9_0_14_cascade_));
    InMux I__7355 (
            .O(N__38366),
            .I(N__38363));
    LocalMux I__7354 (
            .O(N__38363),
            .I(N__38360));
    Span4Mux_h I__7353 (
            .O(N__38360),
            .I(N__38357));
    Odrv4 I__7352 (
            .O(N__38357),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ));
    InMux I__7351 (
            .O(N__38354),
            .I(N__38350));
    InMux I__7350 (
            .O(N__38353),
            .I(N__38347));
    LocalMux I__7349 (
            .O(N__38350),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    LocalMux I__7348 (
            .O(N__38347),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    InMux I__7347 (
            .O(N__38342),
            .I(N__38338));
    CascadeMux I__7346 (
            .O(N__38341),
            .I(N__38335));
    LocalMux I__7345 (
            .O(N__38338),
            .I(N__38331));
    InMux I__7344 (
            .O(N__38335),
            .I(N__38326));
    InMux I__7343 (
            .O(N__38334),
            .I(N__38326));
    Span4Mux_v I__7342 (
            .O(N__38331),
            .I(N__38323));
    LocalMux I__7341 (
            .O(N__38326),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv4 I__7340 (
            .O(N__38323),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    InMux I__7339 (
            .O(N__38318),
            .I(N__38314));
    InMux I__7338 (
            .O(N__38317),
            .I(N__38311));
    LocalMux I__7337 (
            .O(N__38314),
            .I(N__38307));
    LocalMux I__7336 (
            .O(N__38311),
            .I(N__38304));
    InMux I__7335 (
            .O(N__38310),
            .I(N__38301));
    Span4Mux_v I__7334 (
            .O(N__38307),
            .I(N__38298));
    Sp12to4 I__7333 (
            .O(N__38304),
            .I(N__38293));
    LocalMux I__7332 (
            .O(N__38301),
            .I(N__38293));
    Odrv4 I__7331 (
            .O(N__38298),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv12 I__7330 (
            .O(N__38293),
            .I(\current_shift_inst.un4_control_input1_17 ));
    ClkMux I__7329 (
            .O(N__38288),
            .I(N__38282));
    ClkMux I__7328 (
            .O(N__38287),
            .I(N__38282));
    GlobalMux I__7327 (
            .O(N__38282),
            .I(N__38279));
    gio2CtrlBuf I__7326 (
            .O(N__38279),
            .I(delay_hc_input_c_g));
    InMux I__7325 (
            .O(N__38276),
            .I(N__38273));
    LocalMux I__7324 (
            .O(N__38273),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    InMux I__7323 (
            .O(N__38270),
            .I(N__38266));
    InMux I__7322 (
            .O(N__38269),
            .I(N__38263));
    LocalMux I__7321 (
            .O(N__38266),
            .I(N__38259));
    LocalMux I__7320 (
            .O(N__38263),
            .I(N__38256));
    InMux I__7319 (
            .O(N__38262),
            .I(N__38253));
    Span4Mux_v I__7318 (
            .O(N__38259),
            .I(N__38248));
    Span4Mux_v I__7317 (
            .O(N__38256),
            .I(N__38248));
    LocalMux I__7316 (
            .O(N__38253),
            .I(\current_shift_inst.un4_control_input1_9 ));
    Odrv4 I__7315 (
            .O(N__38248),
            .I(\current_shift_inst.un4_control_input1_9 ));
    CascadeMux I__7314 (
            .O(N__38243),
            .I(N__38239));
    InMux I__7313 (
            .O(N__38242),
            .I(N__38233));
    InMux I__7312 (
            .O(N__38239),
            .I(N__38233));
    InMux I__7311 (
            .O(N__38238),
            .I(N__38230));
    LocalMux I__7310 (
            .O(N__38233),
            .I(N__38227));
    LocalMux I__7309 (
            .O(N__38230),
            .I(N__38224));
    Odrv4 I__7308 (
            .O(N__38227),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv12 I__7307 (
            .O(N__38224),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__7306 (
            .O(N__38219),
            .I(N__38216));
    LocalMux I__7305 (
            .O(N__38216),
            .I(N__38211));
    InMux I__7304 (
            .O(N__38215),
            .I(N__38208));
    InMux I__7303 (
            .O(N__38214),
            .I(N__38205));
    Sp12to4 I__7302 (
            .O(N__38211),
            .I(N__38200));
    LocalMux I__7301 (
            .O(N__38208),
            .I(N__38200));
    LocalMux I__7300 (
            .O(N__38205),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv12 I__7299 (
            .O(N__38200),
            .I(\current_shift_inst.un4_control_input1_26 ));
    CascadeMux I__7298 (
            .O(N__38195),
            .I(N__38190));
    InMux I__7297 (
            .O(N__38194),
            .I(N__38187));
    InMux I__7296 (
            .O(N__38193),
            .I(N__38182));
    InMux I__7295 (
            .O(N__38190),
            .I(N__38182));
    LocalMux I__7294 (
            .O(N__38187),
            .I(N__38179));
    LocalMux I__7293 (
            .O(N__38182),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv12 I__7292 (
            .O(N__38179),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__7291 (
            .O(N__38174),
            .I(N__38169));
    InMux I__7290 (
            .O(N__38173),
            .I(N__38166));
    InMux I__7289 (
            .O(N__38172),
            .I(N__38163));
    LocalMux I__7288 (
            .O(N__38169),
            .I(N__38160));
    LocalMux I__7287 (
            .O(N__38166),
            .I(N__38157));
    LocalMux I__7286 (
            .O(N__38163),
            .I(N__38154));
    Odrv4 I__7285 (
            .O(N__38160),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__7284 (
            .O(N__38157),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__7283 (
            .O(N__38154),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__7282 (
            .O(N__38147),
            .I(N__38141));
    InMux I__7281 (
            .O(N__38146),
            .I(N__38141));
    LocalMux I__7280 (
            .O(N__38141),
            .I(N__38137));
    InMux I__7279 (
            .O(N__38140),
            .I(N__38134));
    Sp12to4 I__7278 (
            .O(N__38137),
            .I(N__38129));
    LocalMux I__7277 (
            .O(N__38134),
            .I(N__38129));
    Odrv12 I__7276 (
            .O(N__38129),
            .I(\current_shift_inst.un4_control_input1_2 ));
    CascadeMux I__7275 (
            .O(N__38126),
            .I(N__38121));
    InMux I__7274 (
            .O(N__38125),
            .I(N__38117));
    InMux I__7273 (
            .O(N__38124),
            .I(N__38114));
    InMux I__7272 (
            .O(N__38121),
            .I(N__38111));
    InMux I__7271 (
            .O(N__38120),
            .I(N__38108));
    LocalMux I__7270 (
            .O(N__38117),
            .I(N__38105));
    LocalMux I__7269 (
            .O(N__38114),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__7268 (
            .O(N__38111),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__7267 (
            .O(N__38108),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    Odrv4 I__7266 (
            .O(N__38105),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__7265 (
            .O(N__38096),
            .I(N__38093));
    InMux I__7264 (
            .O(N__38093),
            .I(N__38088));
    InMux I__7263 (
            .O(N__38092),
            .I(N__38085));
    InMux I__7262 (
            .O(N__38091),
            .I(N__38082));
    LocalMux I__7261 (
            .O(N__38088),
            .I(N__38075));
    LocalMux I__7260 (
            .O(N__38085),
            .I(N__38075));
    LocalMux I__7259 (
            .O(N__38082),
            .I(N__38075));
    Odrv12 I__7258 (
            .O(N__38075),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__7257 (
            .O(N__38072),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__7256 (
            .O(N__38069),
            .I(bfn_14_16_0_));
    InMux I__7255 (
            .O(N__38066),
            .I(N__38063));
    LocalMux I__7254 (
            .O(N__38063),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__7253 (
            .O(N__38060),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__7252 (
            .O(N__38057),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__7251 (
            .O(N__38054),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__7250 (
            .O(N__38051),
            .I(N__38048));
    LocalMux I__7249 (
            .O(N__38048),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__7248 (
            .O(N__38045),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__7247 (
            .O(N__38042),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__7246 (
            .O(N__38039),
            .I(N__38034));
    InMux I__7245 (
            .O(N__38038),
            .I(N__38031));
    InMux I__7244 (
            .O(N__38037),
            .I(N__38028));
    LocalMux I__7243 (
            .O(N__38034),
            .I(N__38023));
    LocalMux I__7242 (
            .O(N__38031),
            .I(N__38023));
    LocalMux I__7241 (
            .O(N__38028),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__7240 (
            .O(N__38023),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__7239 (
            .O(N__38018),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__7238 (
            .O(N__38015),
            .I(N__38012));
    LocalMux I__7237 (
            .O(N__38012),
            .I(N__38009));
    Odrv12 I__7236 (
            .O(N__38009),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__7235 (
            .O(N__38006),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__7234 (
            .O(N__38003),
            .I(bfn_14_15_0_));
    CascadeMux I__7233 (
            .O(N__38000),
            .I(N__37996));
    InMux I__7232 (
            .O(N__37999),
            .I(N__37988));
    InMux I__7231 (
            .O(N__37996),
            .I(N__37988));
    InMux I__7230 (
            .O(N__37995),
            .I(N__37988));
    LocalMux I__7229 (
            .O(N__37988),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__7228 (
            .O(N__37985),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__7227 (
            .O(N__37982),
            .I(N__37979));
    LocalMux I__7226 (
            .O(N__37979),
            .I(N__37976));
    Span4Mux_v I__7225 (
            .O(N__37976),
            .I(N__37973));
    Odrv4 I__7224 (
            .O(N__37973),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__7223 (
            .O(N__37970),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__7222 (
            .O(N__37967),
            .I(N__37964));
    LocalMux I__7221 (
            .O(N__37964),
            .I(N__37961));
    Odrv12 I__7220 (
            .O(N__37961),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__7219 (
            .O(N__37958),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__7218 (
            .O(N__37955),
            .I(N__37952));
    LocalMux I__7217 (
            .O(N__37952),
            .I(N__37949));
    Odrv4 I__7216 (
            .O(N__37949),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__7215 (
            .O(N__37946),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__7214 (
            .O(N__37943),
            .I(N__37940));
    LocalMux I__7213 (
            .O(N__37940),
            .I(N__37937));
    Odrv4 I__7212 (
            .O(N__37937),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__7211 (
            .O(N__37934),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__7210 (
            .O(N__37931),
            .I(N__37928));
    LocalMux I__7209 (
            .O(N__37928),
            .I(N__37925));
    Odrv4 I__7208 (
            .O(N__37925),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__7207 (
            .O(N__37922),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__7206 (
            .O(N__37919),
            .I(N__37916));
    LocalMux I__7205 (
            .O(N__37916),
            .I(N__37913));
    Odrv4 I__7204 (
            .O(N__37913),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__7203 (
            .O(N__37910),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__7202 (
            .O(N__37907),
            .I(N__37904));
    LocalMux I__7201 (
            .O(N__37904),
            .I(N__37901));
    Odrv4 I__7200 (
            .O(N__37901),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__7199 (
            .O(N__37898),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__7198 (
            .O(N__37895),
            .I(bfn_14_14_0_));
    InMux I__7197 (
            .O(N__37892),
            .I(N__37889));
    LocalMux I__7196 (
            .O(N__37889),
            .I(N__37886));
    Odrv12 I__7195 (
            .O(N__37886),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__7194 (
            .O(N__37883),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__7193 (
            .O(N__37880),
            .I(N__37877));
    LocalMux I__7192 (
            .O(N__37877),
            .I(N__37874));
    Odrv4 I__7191 (
            .O(N__37874),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__7190 (
            .O(N__37871),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__7189 (
            .O(N__37868),
            .I(N__37865));
    LocalMux I__7188 (
            .O(N__37865),
            .I(N__37862));
    Odrv4 I__7187 (
            .O(N__37862),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__7186 (
            .O(N__37859),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__7185 (
            .O(N__37856),
            .I(N__37853));
    LocalMux I__7184 (
            .O(N__37853),
            .I(N__37850));
    Span4Mux_v I__7183 (
            .O(N__37850),
            .I(N__37847));
    Odrv4 I__7182 (
            .O(N__37847),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__7181 (
            .O(N__37844),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__7180 (
            .O(N__37841),
            .I(N__37838));
    LocalMux I__7179 (
            .O(N__37838),
            .I(N__37835));
    Odrv12 I__7178 (
            .O(N__37835),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__7177 (
            .O(N__37832),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__7176 (
            .O(N__37829),
            .I(N__37826));
    LocalMux I__7175 (
            .O(N__37826),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__7174 (
            .O(N__37823),
            .I(N__37817));
    InMux I__7173 (
            .O(N__37822),
            .I(N__37814));
    InMux I__7172 (
            .O(N__37821),
            .I(N__37811));
    InMux I__7171 (
            .O(N__37820),
            .I(N__37808));
    InMux I__7170 (
            .O(N__37817),
            .I(N__37805));
    LocalMux I__7169 (
            .O(N__37814),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__7168 (
            .O(N__37811),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__7167 (
            .O(N__37808),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__7166 (
            .O(N__37805),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__7165 (
            .O(N__37796),
            .I(N__37793));
    LocalMux I__7164 (
            .O(N__37793),
            .I(N__37790));
    Odrv4 I__7163 (
            .O(N__37790),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__7162 (
            .O(N__37787),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__7161 (
            .O(N__37784),
            .I(N__37781));
    LocalMux I__7160 (
            .O(N__37781),
            .I(N__37778));
    Odrv4 I__7159 (
            .O(N__37778),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__7158 (
            .O(N__37775),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__7157 (
            .O(N__37772),
            .I(N__37769));
    LocalMux I__7156 (
            .O(N__37769),
            .I(N__37766));
    Odrv4 I__7155 (
            .O(N__37766),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__7154 (
            .O(N__37763),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__7153 (
            .O(N__37760),
            .I(N__37757));
    LocalMux I__7152 (
            .O(N__37757),
            .I(N__37754));
    Odrv4 I__7151 (
            .O(N__37754),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__7150 (
            .O(N__37751),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__7149 (
            .O(N__37748),
            .I(N__37745));
    LocalMux I__7148 (
            .O(N__37745),
            .I(N__37742));
    Odrv4 I__7147 (
            .O(N__37742),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__7146 (
            .O(N__37739),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__7145 (
            .O(N__37736),
            .I(N__37732));
    InMux I__7144 (
            .O(N__37735),
            .I(N__37726));
    LocalMux I__7143 (
            .O(N__37732),
            .I(N__37723));
    InMux I__7142 (
            .O(N__37731),
            .I(N__37720));
    CascadeMux I__7141 (
            .O(N__37730),
            .I(N__37716));
    InMux I__7140 (
            .O(N__37729),
            .I(N__37713));
    LocalMux I__7139 (
            .O(N__37726),
            .I(N__37710));
    Span4Mux_v I__7138 (
            .O(N__37723),
            .I(N__37707));
    LocalMux I__7137 (
            .O(N__37720),
            .I(N__37704));
    InMux I__7136 (
            .O(N__37719),
            .I(N__37701));
    InMux I__7135 (
            .O(N__37716),
            .I(N__37698));
    LocalMux I__7134 (
            .O(N__37713),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__7133 (
            .O(N__37710),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__7132 (
            .O(N__37707),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv12 I__7131 (
            .O(N__37704),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    LocalMux I__7130 (
            .O(N__37701),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    LocalMux I__7129 (
            .O(N__37698),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__7128 (
            .O(N__37685),
            .I(N__37682));
    LocalMux I__7127 (
            .O(N__37682),
            .I(N__37677));
    CascadeMux I__7126 (
            .O(N__37681),
            .I(N__37674));
    InMux I__7125 (
            .O(N__37680),
            .I(N__37671));
    Span4Mux_v I__7124 (
            .O(N__37677),
            .I(N__37668));
    InMux I__7123 (
            .O(N__37674),
            .I(N__37665));
    LocalMux I__7122 (
            .O(N__37671),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ));
    Odrv4 I__7121 (
            .O(N__37668),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ));
    LocalMux I__7120 (
            .O(N__37665),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ));
    InMux I__7119 (
            .O(N__37658),
            .I(N__37655));
    LocalMux I__7118 (
            .O(N__37655),
            .I(N__37652));
    Odrv12 I__7117 (
            .O(N__37652),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ));
    CEMux I__7116 (
            .O(N__37649),
            .I(N__37644));
    CEMux I__7115 (
            .O(N__37648),
            .I(N__37639));
    CEMux I__7114 (
            .O(N__37647),
            .I(N__37636));
    LocalMux I__7113 (
            .O(N__37644),
            .I(N__37632));
    CEMux I__7112 (
            .O(N__37643),
            .I(N__37629));
    CEMux I__7111 (
            .O(N__37642),
            .I(N__37626));
    LocalMux I__7110 (
            .O(N__37639),
            .I(N__37623));
    LocalMux I__7109 (
            .O(N__37636),
            .I(N__37619));
    CEMux I__7108 (
            .O(N__37635),
            .I(N__37616));
    Span4Mux_h I__7107 (
            .O(N__37632),
            .I(N__37613));
    LocalMux I__7106 (
            .O(N__37629),
            .I(N__37610));
    LocalMux I__7105 (
            .O(N__37626),
            .I(N__37607));
    Span4Mux_h I__7104 (
            .O(N__37623),
            .I(N__37604));
    CEMux I__7103 (
            .O(N__37622),
            .I(N__37601));
    Span4Mux_v I__7102 (
            .O(N__37619),
            .I(N__37595));
    LocalMux I__7101 (
            .O(N__37616),
            .I(N__37595));
    Span4Mux_v I__7100 (
            .O(N__37613),
            .I(N__37590));
    Span4Mux_h I__7099 (
            .O(N__37610),
            .I(N__37590));
    Span4Mux_v I__7098 (
            .O(N__37607),
            .I(N__37587));
    Sp12to4 I__7097 (
            .O(N__37604),
            .I(N__37582));
    LocalMux I__7096 (
            .O(N__37601),
            .I(N__37582));
    CEMux I__7095 (
            .O(N__37600),
            .I(N__37579));
    Odrv4 I__7094 (
            .O(N__37595),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__7093 (
            .O(N__37590),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__7092 (
            .O(N__37587),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv12 I__7091 (
            .O(N__37582),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    LocalMux I__7090 (
            .O(N__37579),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    CascadeMux I__7089 (
            .O(N__37568),
            .I(elapsed_time_ns_1_RNI46CN9_0_17_cascade_));
    InMux I__7088 (
            .O(N__37565),
            .I(N__37562));
    LocalMux I__7087 (
            .O(N__37562),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ));
    InMux I__7086 (
            .O(N__37559),
            .I(N__37556));
    LocalMux I__7085 (
            .O(N__37556),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ));
    InMux I__7084 (
            .O(N__37553),
            .I(N__37550));
    LocalMux I__7083 (
            .O(N__37550),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ));
    CascadeMux I__7082 (
            .O(N__37547),
            .I(elapsed_time_ns_1_RNIL73T9_0_9_cascade_));
    InMux I__7081 (
            .O(N__37544),
            .I(N__37541));
    LocalMux I__7080 (
            .O(N__37541),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ));
    InMux I__7079 (
            .O(N__37538),
            .I(N__37535));
    LocalMux I__7078 (
            .O(N__37535),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    CascadeMux I__7077 (
            .O(N__37532),
            .I(elapsed_time_ns_1_RNI14DN9_0_23_cascade_));
    InMux I__7076 (
            .O(N__37529),
            .I(N__37526));
    LocalMux I__7075 (
            .O(N__37526),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ));
    InMux I__7074 (
            .O(N__37523),
            .I(N__37520));
    LocalMux I__7073 (
            .O(N__37520),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ));
    InMux I__7072 (
            .O(N__37517),
            .I(N__37514));
    LocalMux I__7071 (
            .O(N__37514),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    CascadeMux I__7070 (
            .O(N__37511),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21_cascade_));
    InMux I__7069 (
            .O(N__37508),
            .I(N__37505));
    LocalMux I__7068 (
            .O(N__37505),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ));
    InMux I__7067 (
            .O(N__37502),
            .I(N__37499));
    LocalMux I__7066 (
            .O(N__37499),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ));
    InMux I__7065 (
            .O(N__37496),
            .I(N__37493));
    LocalMux I__7064 (
            .O(N__37493),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    InMux I__7063 (
            .O(N__37490),
            .I(N__37487));
    LocalMux I__7062 (
            .O(N__37487),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ));
    InMux I__7061 (
            .O(N__37484),
            .I(N__37480));
    InMux I__7060 (
            .O(N__37483),
            .I(N__37477));
    LocalMux I__7059 (
            .O(N__37480),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    LocalMux I__7058 (
            .O(N__37477),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__7057 (
            .O(N__37472),
            .I(N__37468));
    InMux I__7056 (
            .O(N__37471),
            .I(N__37465));
    LocalMux I__7055 (
            .O(N__37468),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    LocalMux I__7054 (
            .O(N__37465),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__7053 (
            .O(N__37460),
            .I(N__37457));
    LocalMux I__7052 (
            .O(N__37457),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    CascadeMux I__7051 (
            .O(N__37454),
            .I(elapsed_time_ns_1_RNI47DN9_0_26_cascade_));
    CascadeMux I__7050 (
            .O(N__37451),
            .I(N__37448));
    InMux I__7049 (
            .O(N__37448),
            .I(N__37445));
    LocalMux I__7048 (
            .O(N__37445),
            .I(N__37442));
    Odrv4 I__7047 (
            .O(N__37442),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ));
    InMux I__7046 (
            .O(N__37439),
            .I(N__37435));
    InMux I__7045 (
            .O(N__37438),
            .I(N__37432));
    LocalMux I__7044 (
            .O(N__37435),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__7043 (
            .O(N__37432),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    InMux I__7042 (
            .O(N__37427),
            .I(N__37424));
    LocalMux I__7041 (
            .O(N__37424),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ));
    InMux I__7040 (
            .O(N__37421),
            .I(N__37418));
    LocalMux I__7039 (
            .O(N__37418),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ));
    InMux I__7038 (
            .O(N__37415),
            .I(N__37412));
    LocalMux I__7037 (
            .O(N__37412),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ));
    InMux I__7036 (
            .O(N__37409),
            .I(N__37406));
    LocalMux I__7035 (
            .O(N__37406),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    InMux I__7034 (
            .O(N__37403),
            .I(N__37400));
    LocalMux I__7033 (
            .O(N__37400),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    CascadeMux I__7032 (
            .O(N__37397),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11_cascade_));
    CascadeMux I__7031 (
            .O(N__37394),
            .I(N__37391));
    InMux I__7030 (
            .O(N__37391),
            .I(N__37388));
    LocalMux I__7029 (
            .O(N__37388),
            .I(N__37385));
    Odrv4 I__7028 (
            .O(N__37385),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ));
    InMux I__7027 (
            .O(N__37382),
            .I(N__37379));
    LocalMux I__7026 (
            .O(N__37379),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    CascadeMux I__7025 (
            .O(N__37376),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_));
    InMux I__7024 (
            .O(N__37373),
            .I(N__37370));
    LocalMux I__7023 (
            .O(N__37370),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ));
    InMux I__7022 (
            .O(N__37367),
            .I(N__37364));
    LocalMux I__7021 (
            .O(N__37364),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    CascadeMux I__7020 (
            .O(N__37361),
            .I(elapsed_time_ns_1_RNIK63T9_0_8_cascade_));
    InMux I__7019 (
            .O(N__37358),
            .I(N__37355));
    LocalMux I__7018 (
            .O(N__37355),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ));
    InMux I__7017 (
            .O(N__37352),
            .I(N__37348));
    InMux I__7016 (
            .O(N__37351),
            .I(N__37345));
    LocalMux I__7015 (
            .O(N__37348),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__7014 (
            .O(N__37345),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    InMux I__7013 (
            .O(N__37340),
            .I(N__37337));
    LocalMux I__7012 (
            .O(N__37337),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ));
    InMux I__7011 (
            .O(N__37334),
            .I(N__37331));
    LocalMux I__7010 (
            .O(N__37331),
            .I(N__37328));
    Span12Mux_s6_h I__7009 (
            .O(N__37328),
            .I(N__37325));
    Odrv12 I__7008 (
            .O(N__37325),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ));
    InMux I__7007 (
            .O(N__37322),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    InMux I__7006 (
            .O(N__37319),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    InMux I__7005 (
            .O(N__37316),
            .I(N__37313));
    LocalMux I__7004 (
            .O(N__37313),
            .I(N__37310));
    Span12Mux_s5_h I__7003 (
            .O(N__37310),
            .I(N__37307));
    Odrv12 I__7002 (
            .O(N__37307),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO ));
    InMux I__7001 (
            .O(N__37304),
            .I(N__37301));
    LocalMux I__7000 (
            .O(N__37301),
            .I(N__37297));
    InMux I__6999 (
            .O(N__37300),
            .I(N__37294));
    Span4Mux_v I__6998 (
            .O(N__37297),
            .I(N__37288));
    LocalMux I__6997 (
            .O(N__37294),
            .I(N__37288));
    InMux I__6996 (
            .O(N__37293),
            .I(N__37284));
    Span4Mux_v I__6995 (
            .O(N__37288),
            .I(N__37281));
    CascadeMux I__6994 (
            .O(N__37287),
            .I(N__37278));
    LocalMux I__6993 (
            .O(N__37284),
            .I(N__37273));
    Span4Mux_h I__6992 (
            .O(N__37281),
            .I(N__37270));
    InMux I__6991 (
            .O(N__37278),
            .I(N__37263));
    InMux I__6990 (
            .O(N__37277),
            .I(N__37263));
    InMux I__6989 (
            .O(N__37276),
            .I(N__37263));
    Span12Mux_v I__6988 (
            .O(N__37273),
            .I(N__37260));
    Span4Mux_v I__6987 (
            .O(N__37270),
            .I(N__37257));
    LocalMux I__6986 (
            .O(N__37263),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__6985 (
            .O(N__37260),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__6984 (
            .O(N__37257),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__6983 (
            .O(N__37250),
            .I(N__37244));
    InMux I__6982 (
            .O(N__37249),
            .I(N__37244));
    LocalMux I__6981 (
            .O(N__37244),
            .I(N__37239));
    InMux I__6980 (
            .O(N__37243),
            .I(N__37235));
    InMux I__6979 (
            .O(N__37242),
            .I(N__37232));
    Span12Mux_h I__6978 (
            .O(N__37239),
            .I(N__37228));
    InMux I__6977 (
            .O(N__37238),
            .I(N__37225));
    LocalMux I__6976 (
            .O(N__37235),
            .I(N__37222));
    LocalMux I__6975 (
            .O(N__37232),
            .I(N__37219));
    InMux I__6974 (
            .O(N__37231),
            .I(N__37216));
    Span12Mux_v I__6973 (
            .O(N__37228),
            .I(N__37211));
    LocalMux I__6972 (
            .O(N__37225),
            .I(N__37211));
    Span4Mux_v I__6971 (
            .O(N__37222),
            .I(N__37206));
    Span4Mux_v I__6970 (
            .O(N__37219),
            .I(N__37206));
    LocalMux I__6969 (
            .O(N__37216),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv12 I__6968 (
            .O(N__37211),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__6967 (
            .O(N__37206),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__6966 (
            .O(N__37199),
            .I(N__37195));
    InMux I__6965 (
            .O(N__37198),
            .I(N__37192));
    LocalMux I__6964 (
            .O(N__37195),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    LocalMux I__6963 (
            .O(N__37192),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__6962 (
            .O(N__37187),
            .I(N__37184));
    LocalMux I__6961 (
            .O(N__37184),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    CascadeMux I__6960 (
            .O(N__37181),
            .I(elapsed_time_ns_1_RNITUBN9_0_10_cascade_));
    InMux I__6959 (
            .O(N__37178),
            .I(N__37175));
    LocalMux I__6958 (
            .O(N__37175),
            .I(N__37172));
    Odrv4 I__6957 (
            .O(N__37172),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ));
    InMux I__6956 (
            .O(N__37169),
            .I(N__37166));
    LocalMux I__6955 (
            .O(N__37166),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ));
    InMux I__6954 (
            .O(N__37163),
            .I(N__37160));
    LocalMux I__6953 (
            .O(N__37160),
            .I(N__37157));
    Span4Mux_v I__6952 (
            .O(N__37157),
            .I(N__37154));
    Span4Mux_h I__6951 (
            .O(N__37154),
            .I(N__37151));
    Span4Mux_h I__6950 (
            .O(N__37151),
            .I(N__37148));
    Span4Mux_h I__6949 (
            .O(N__37148),
            .I(N__37145));
    Odrv4 I__6948 (
            .O(N__37145),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    InMux I__6947 (
            .O(N__37142),
            .I(N__37139));
    LocalMux I__6946 (
            .O(N__37139),
            .I(N__37136));
    Span12Mux_s5_h I__6945 (
            .O(N__37136),
            .I(N__37133));
    Odrv12 I__6944 (
            .O(N__37133),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ));
    InMux I__6943 (
            .O(N__37130),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    CascadeMux I__6942 (
            .O(N__37127),
            .I(N__37124));
    InMux I__6941 (
            .O(N__37124),
            .I(N__37121));
    LocalMux I__6940 (
            .O(N__37121),
            .I(N__37118));
    Span4Mux_v I__6939 (
            .O(N__37118),
            .I(N__37115));
    Span4Mux_v I__6938 (
            .O(N__37115),
            .I(N__37112));
    Sp12to4 I__6937 (
            .O(N__37112),
            .I(N__37109));
    Odrv12 I__6936 (
            .O(N__37109),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    InMux I__6935 (
            .O(N__37106),
            .I(N__37103));
    LocalMux I__6934 (
            .O(N__37103),
            .I(N__37100));
    Span12Mux_s4_h I__6933 (
            .O(N__37100),
            .I(N__37097));
    Odrv12 I__6932 (
            .O(N__37097),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ));
    InMux I__6931 (
            .O(N__37094),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__6930 (
            .O(N__37091),
            .I(N__37088));
    LocalMux I__6929 (
            .O(N__37088),
            .I(N__37085));
    Span12Mux_h I__6928 (
            .O(N__37085),
            .I(N__37082));
    Span12Mux_h I__6927 (
            .O(N__37082),
            .I(N__37079));
    Odrv12 I__6926 (
            .O(N__37079),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    InMux I__6925 (
            .O(N__37076),
            .I(N__37073));
    LocalMux I__6924 (
            .O(N__37073),
            .I(N__37070));
    Span12Mux_s3_h I__6923 (
            .O(N__37070),
            .I(N__37067));
    Odrv12 I__6922 (
            .O(N__37067),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ));
    InMux I__6921 (
            .O(N__37064),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    CascadeMux I__6920 (
            .O(N__37061),
            .I(N__37058));
    InMux I__6919 (
            .O(N__37058),
            .I(N__37055));
    LocalMux I__6918 (
            .O(N__37055),
            .I(N__37052));
    Span4Mux_v I__6917 (
            .O(N__37052),
            .I(N__37049));
    Span4Mux_h I__6916 (
            .O(N__37049),
            .I(N__37046));
    Span4Mux_h I__6915 (
            .O(N__37046),
            .I(N__37043));
    Span4Mux_h I__6914 (
            .O(N__37043),
            .I(N__37040));
    Odrv4 I__6913 (
            .O(N__37040),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    InMux I__6912 (
            .O(N__37037),
            .I(N__37034));
    LocalMux I__6911 (
            .O(N__37034),
            .I(N__37031));
    Span12Mux_s2_h I__6910 (
            .O(N__37031),
            .I(N__37028));
    Odrv12 I__6909 (
            .O(N__37028),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ));
    InMux I__6908 (
            .O(N__37025),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    CascadeMux I__6907 (
            .O(N__37022),
            .I(N__37019));
    InMux I__6906 (
            .O(N__37019),
            .I(N__37016));
    LocalMux I__6905 (
            .O(N__37016),
            .I(N__37013));
    Span4Mux_v I__6904 (
            .O(N__37013),
            .I(N__37010));
    Sp12to4 I__6903 (
            .O(N__37010),
            .I(N__37007));
    Span12Mux_h I__6902 (
            .O(N__37007),
            .I(N__37004));
    Odrv12 I__6901 (
            .O(N__37004),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    InMux I__6900 (
            .O(N__37001),
            .I(N__36998));
    LocalMux I__6899 (
            .O(N__36998),
            .I(N__36995));
    Span12Mux_s9_h I__6898 (
            .O(N__36995),
            .I(N__36992));
    Odrv12 I__6897 (
            .O(N__36992),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ));
    InMux I__6896 (
            .O(N__36989),
            .I(bfn_13_22_0_));
    InMux I__6895 (
            .O(N__36986),
            .I(N__36983));
    LocalMux I__6894 (
            .O(N__36983),
            .I(N__36980));
    Span4Mux_v I__6893 (
            .O(N__36980),
            .I(N__36977));
    Sp12to4 I__6892 (
            .O(N__36977),
            .I(N__36974));
    Span12Mux_h I__6891 (
            .O(N__36974),
            .I(N__36971));
    Odrv12 I__6890 (
            .O(N__36971),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    InMux I__6889 (
            .O(N__36968),
            .I(N__36965));
    LocalMux I__6888 (
            .O(N__36965),
            .I(N__36962));
    Span12Mux_s8_h I__6887 (
            .O(N__36962),
            .I(N__36959));
    Odrv12 I__6886 (
            .O(N__36959),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ));
    InMux I__6885 (
            .O(N__36956),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    InMux I__6884 (
            .O(N__36953),
            .I(N__36950));
    LocalMux I__6883 (
            .O(N__36950),
            .I(N__36947));
    Span4Mux_h I__6882 (
            .O(N__36947),
            .I(N__36944));
    Span4Mux_h I__6881 (
            .O(N__36944),
            .I(N__36941));
    Sp12to4 I__6880 (
            .O(N__36941),
            .I(N__36938));
    Span12Mux_v I__6879 (
            .O(N__36938),
            .I(N__36935));
    Odrv12 I__6878 (
            .O(N__36935),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__6877 (
            .O(N__36932),
            .I(N__36929));
    LocalMux I__6876 (
            .O(N__36929),
            .I(N__36926));
    Span12Mux_s7_h I__6875 (
            .O(N__36926),
            .I(N__36923));
    Odrv12 I__6874 (
            .O(N__36923),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ));
    InMux I__6873 (
            .O(N__36920),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    InMux I__6872 (
            .O(N__36917),
            .I(N__36914));
    LocalMux I__6871 (
            .O(N__36914),
            .I(N__36911));
    Span4Mux_v I__6870 (
            .O(N__36911),
            .I(N__36908));
    Sp12to4 I__6869 (
            .O(N__36908),
            .I(N__36905));
    Span12Mux_h I__6868 (
            .O(N__36905),
            .I(N__36902));
    Odrv12 I__6867 (
            .O(N__36902),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    CascadeMux I__6866 (
            .O(N__36899),
            .I(N__36893));
    CascadeMux I__6865 (
            .O(N__36898),
            .I(N__36890));
    CascadeMux I__6864 (
            .O(N__36897),
            .I(N__36887));
    CascadeMux I__6863 (
            .O(N__36896),
            .I(N__36881));
    InMux I__6862 (
            .O(N__36893),
            .I(N__36878));
    InMux I__6861 (
            .O(N__36890),
            .I(N__36871));
    InMux I__6860 (
            .O(N__36887),
            .I(N__36871));
    InMux I__6859 (
            .O(N__36886),
            .I(N__36871));
    CascadeMux I__6858 (
            .O(N__36885),
            .I(N__36867));
    CascadeMux I__6857 (
            .O(N__36884),
            .I(N__36863));
    InMux I__6856 (
            .O(N__36881),
            .I(N__36860));
    LocalMux I__6855 (
            .O(N__36878),
            .I(N__36857));
    LocalMux I__6854 (
            .O(N__36871),
            .I(N__36854));
    InMux I__6853 (
            .O(N__36870),
            .I(N__36845));
    InMux I__6852 (
            .O(N__36867),
            .I(N__36845));
    InMux I__6851 (
            .O(N__36866),
            .I(N__36845));
    InMux I__6850 (
            .O(N__36863),
            .I(N__36845));
    LocalMux I__6849 (
            .O(N__36860),
            .I(N__36842));
    Span4Mux_v I__6848 (
            .O(N__36857),
            .I(N__36835));
    Span4Mux_v I__6847 (
            .O(N__36854),
            .I(N__36835));
    LocalMux I__6846 (
            .O(N__36845),
            .I(N__36835));
    Span12Mux_s10_v I__6845 (
            .O(N__36842),
            .I(N__36832));
    Span4Mux_v I__6844 (
            .O(N__36835),
            .I(N__36829));
    Span12Mux_h I__6843 (
            .O(N__36832),
            .I(N__36826));
    Span4Mux_h I__6842 (
            .O(N__36829),
            .I(N__36823));
    Span12Mux_h I__6841 (
            .O(N__36826),
            .I(N__36820));
    Span4Mux_h I__6840 (
            .O(N__36823),
            .I(N__36817));
    Odrv12 I__6839 (
            .O(N__36820),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    Odrv4 I__6838 (
            .O(N__36817),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__6837 (
            .O(N__36812),
            .I(N__36809));
    LocalMux I__6836 (
            .O(N__36809),
            .I(N__36806));
    Span4Mux_v I__6835 (
            .O(N__36806),
            .I(N__36803));
    Span4Mux_h I__6834 (
            .O(N__36803),
            .I(N__36800));
    Span4Mux_h I__6833 (
            .O(N__36800),
            .I(N__36797));
    Span4Mux_h I__6832 (
            .O(N__36797),
            .I(N__36794));
    Odrv4 I__6831 (
            .O(N__36794),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__6830 (
            .O(N__36791),
            .I(N__36788));
    InMux I__6829 (
            .O(N__36788),
            .I(N__36785));
    LocalMux I__6828 (
            .O(N__36785),
            .I(N__36782));
    Sp12to4 I__6827 (
            .O(N__36782),
            .I(N__36779));
    Span12Mux_v I__6826 (
            .O(N__36779),
            .I(N__36776));
    Odrv12 I__6825 (
            .O(N__36776),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    CascadeMux I__6824 (
            .O(N__36773),
            .I(N__36770));
    InMux I__6823 (
            .O(N__36770),
            .I(N__36767));
    LocalMux I__6822 (
            .O(N__36767),
            .I(N__36764));
    Span12Mux_s9_h I__6821 (
            .O(N__36764),
            .I(N__36761));
    Odrv12 I__6820 (
            .O(N__36761),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_8 ));
    InMux I__6819 (
            .O(N__36758),
            .I(N__36755));
    LocalMux I__6818 (
            .O(N__36755),
            .I(N__36752));
    Span4Mux_v I__6817 (
            .O(N__36752),
            .I(N__36749));
    Sp12to4 I__6816 (
            .O(N__36749),
            .I(N__36746));
    Span12Mux_h I__6815 (
            .O(N__36746),
            .I(N__36743));
    Odrv12 I__6814 (
            .O(N__36743),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__6813 (
            .O(N__36740),
            .I(N__36737));
    InMux I__6812 (
            .O(N__36737),
            .I(N__36734));
    LocalMux I__6811 (
            .O(N__36734),
            .I(N__36731));
    Span12Mux_v I__6810 (
            .O(N__36731),
            .I(N__36728));
    Span12Mux_h I__6809 (
            .O(N__36728),
            .I(N__36725));
    Odrv12 I__6808 (
            .O(N__36725),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    CascadeMux I__6807 (
            .O(N__36722),
            .I(N__36719));
    InMux I__6806 (
            .O(N__36719),
            .I(N__36716));
    LocalMux I__6805 (
            .O(N__36716),
            .I(N__36713));
    Span12Mux_s8_h I__6804 (
            .O(N__36713),
            .I(N__36710));
    Odrv12 I__6803 (
            .O(N__36710),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ));
    InMux I__6802 (
            .O(N__36707),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__6801 (
            .O(N__36704),
            .I(N__36701));
    LocalMux I__6800 (
            .O(N__36701),
            .I(N__36698));
    Span4Mux_h I__6799 (
            .O(N__36698),
            .I(N__36695));
    Span4Mux_h I__6798 (
            .O(N__36695),
            .I(N__36692));
    Sp12to4 I__6797 (
            .O(N__36692),
            .I(N__36689));
    Span12Mux_v I__6796 (
            .O(N__36689),
            .I(N__36686));
    Odrv12 I__6795 (
            .O(N__36686),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__6794 (
            .O(N__36683),
            .I(N__36680));
    InMux I__6793 (
            .O(N__36680),
            .I(N__36677));
    LocalMux I__6792 (
            .O(N__36677),
            .I(N__36674));
    Span12Mux_v I__6791 (
            .O(N__36674),
            .I(N__36671));
    Span12Mux_h I__6790 (
            .O(N__36671),
            .I(N__36668));
    Odrv12 I__6789 (
            .O(N__36668),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    CascadeMux I__6788 (
            .O(N__36665),
            .I(N__36662));
    InMux I__6787 (
            .O(N__36662),
            .I(N__36659));
    LocalMux I__6786 (
            .O(N__36659),
            .I(N__36656));
    Span12Mux_s7_h I__6785 (
            .O(N__36656),
            .I(N__36653));
    Odrv12 I__6784 (
            .O(N__36653),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ));
    InMux I__6783 (
            .O(N__36650),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__6782 (
            .O(N__36647),
            .I(N__36644));
    LocalMux I__6781 (
            .O(N__36644),
            .I(N__36641));
    Span4Mux_v I__6780 (
            .O(N__36641),
            .I(N__36638));
    Sp12to4 I__6779 (
            .O(N__36638),
            .I(N__36635));
    Span12Mux_h I__6778 (
            .O(N__36635),
            .I(N__36632));
    Odrv12 I__6777 (
            .O(N__36632),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__6776 (
            .O(N__36629),
            .I(N__36626));
    InMux I__6775 (
            .O(N__36626),
            .I(N__36623));
    LocalMux I__6774 (
            .O(N__36623),
            .I(N__36620));
    Span4Mux_v I__6773 (
            .O(N__36620),
            .I(N__36617));
    Span4Mux_h I__6772 (
            .O(N__36617),
            .I(N__36614));
    Span4Mux_h I__6771 (
            .O(N__36614),
            .I(N__36611));
    Odrv4 I__6770 (
            .O(N__36611),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    CascadeMux I__6769 (
            .O(N__36608),
            .I(N__36605));
    InMux I__6768 (
            .O(N__36605),
            .I(N__36602));
    LocalMux I__6767 (
            .O(N__36602),
            .I(N__36599));
    Span12Mux_s6_h I__6766 (
            .O(N__36599),
            .I(N__36596));
    Odrv12 I__6765 (
            .O(N__36596),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ));
    InMux I__6764 (
            .O(N__36593),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__6763 (
            .O(N__36590),
            .I(N__36584));
    InMux I__6762 (
            .O(N__36589),
            .I(N__36584));
    LocalMux I__6761 (
            .O(N__36584),
            .I(N__36579));
    InMux I__6760 (
            .O(N__36583),
            .I(N__36576));
    InMux I__6759 (
            .O(N__36582),
            .I(N__36573));
    Odrv4 I__6758 (
            .O(N__36579),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6757 (
            .O(N__36576),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6756 (
            .O(N__36573),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__6755 (
            .O(N__36566),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__6754 (
            .O(N__36563),
            .I(N__36560));
    LocalMux I__6753 (
            .O(N__36560),
            .I(\current_shift_inst.un4_control_input1_1 ));
    InMux I__6752 (
            .O(N__36557),
            .I(N__36553));
    InMux I__6751 (
            .O(N__36556),
            .I(N__36550));
    LocalMux I__6750 (
            .O(N__36553),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ));
    LocalMux I__6749 (
            .O(N__36550),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ));
    InMux I__6748 (
            .O(N__36545),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ));
    InMux I__6747 (
            .O(N__36542),
            .I(N__36538));
    InMux I__6746 (
            .O(N__36541),
            .I(N__36535));
    LocalMux I__6745 (
            .O(N__36538),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ));
    LocalMux I__6744 (
            .O(N__36535),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ));
    InMux I__6743 (
            .O(N__36530),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ));
    InMux I__6742 (
            .O(N__36527),
            .I(N__36523));
    InMux I__6741 (
            .O(N__36526),
            .I(N__36520));
    LocalMux I__6740 (
            .O(N__36523),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ));
    LocalMux I__6739 (
            .O(N__36520),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ));
    InMux I__6738 (
            .O(N__36515),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ));
    InMux I__6737 (
            .O(N__36512),
            .I(N__36508));
    InMux I__6736 (
            .O(N__36511),
            .I(N__36505));
    LocalMux I__6735 (
            .O(N__36508),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ));
    LocalMux I__6734 (
            .O(N__36505),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ));
    InMux I__6733 (
            .O(N__36500),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ));
    InMux I__6732 (
            .O(N__36497),
            .I(N__36494));
    LocalMux I__6731 (
            .O(N__36494),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ));
    InMux I__6730 (
            .O(N__36491),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ));
    InMux I__6729 (
            .O(N__36488),
            .I(N__36485));
    LocalMux I__6728 (
            .O(N__36485),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ));
    InMux I__6727 (
            .O(N__36482),
            .I(N__36479));
    LocalMux I__6726 (
            .O(N__36479),
            .I(N__36475));
    InMux I__6725 (
            .O(N__36478),
            .I(N__36472));
    Odrv4 I__6724 (
            .O(N__36475),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_28));
    LocalMux I__6723 (
            .O(N__36472),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_28));
    InMux I__6722 (
            .O(N__36467),
            .I(N__36464));
    LocalMux I__6721 (
            .O(N__36464),
            .I(N__36461));
    Span4Mux_h I__6720 (
            .O(N__36461),
            .I(N__36457));
    InMux I__6719 (
            .O(N__36460),
            .I(N__36453));
    Span4Mux_v I__6718 (
            .O(N__36457),
            .I(N__36450));
    InMux I__6717 (
            .O(N__36456),
            .I(N__36447));
    LocalMux I__6716 (
            .O(N__36453),
            .I(N__36444));
    Span4Mux_v I__6715 (
            .O(N__36450),
            .I(N__36441));
    LocalMux I__6714 (
            .O(N__36447),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ));
    Odrv12 I__6713 (
            .O(N__36444),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ));
    Odrv4 I__6712 (
            .O(N__36441),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ));
    InMux I__6711 (
            .O(N__36434),
            .I(N__36431));
    LocalMux I__6710 (
            .O(N__36431),
            .I(N__36426));
    InMux I__6709 (
            .O(N__36430),
            .I(N__36423));
    InMux I__6708 (
            .O(N__36429),
            .I(N__36420));
    Span12Mux_v I__6707 (
            .O(N__36426),
            .I(N__36417));
    LocalMux I__6706 (
            .O(N__36423),
            .I(N__36414));
    LocalMux I__6705 (
            .O(N__36420),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ));
    Odrv12 I__6704 (
            .O(N__36417),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ));
    Odrv12 I__6703 (
            .O(N__36414),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ));
    InMux I__6702 (
            .O(N__36407),
            .I(N__36398));
    InMux I__6701 (
            .O(N__36406),
            .I(N__36398));
    InMux I__6700 (
            .O(N__36405),
            .I(N__36398));
    LocalMux I__6699 (
            .O(N__36398),
            .I(N__36394));
    InMux I__6698 (
            .O(N__36397),
            .I(N__36391));
    Span4Mux_v I__6697 (
            .O(N__36394),
            .I(N__36388));
    LocalMux I__6696 (
            .O(N__36391),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ));
    Odrv4 I__6695 (
            .O(N__36388),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ));
    CascadeMux I__6694 (
            .O(N__36383),
            .I(N__36380));
    InMux I__6693 (
            .O(N__36380),
            .I(N__36377));
    LocalMux I__6692 (
            .O(N__36377),
            .I(N__36374));
    Span4Mux_h I__6691 (
            .O(N__36374),
            .I(N__36371));
    Odrv4 I__6690 (
            .O(N__36371),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt30 ));
    InMux I__6689 (
            .O(N__36368),
            .I(N__36364));
    InMux I__6688 (
            .O(N__36367),
            .I(N__36361));
    LocalMux I__6687 (
            .O(N__36364),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ));
    LocalMux I__6686 (
            .O(N__36361),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ));
    InMux I__6685 (
            .O(N__36356),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ));
    InMux I__6684 (
            .O(N__36353),
            .I(N__36349));
    InMux I__6683 (
            .O(N__36352),
            .I(N__36346));
    LocalMux I__6682 (
            .O(N__36349),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ));
    LocalMux I__6681 (
            .O(N__36346),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ));
    InMux I__6680 (
            .O(N__36341),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ));
    InMux I__6679 (
            .O(N__36338),
            .I(N__36334));
    InMux I__6678 (
            .O(N__36337),
            .I(N__36331));
    LocalMux I__6677 (
            .O(N__36334),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ));
    LocalMux I__6676 (
            .O(N__36331),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ));
    InMux I__6675 (
            .O(N__36326),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ));
    InMux I__6674 (
            .O(N__36323),
            .I(N__36320));
    LocalMux I__6673 (
            .O(N__36320),
            .I(N__36317));
    Odrv4 I__6672 (
            .O(N__36317),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ));
    InMux I__6671 (
            .O(N__36314),
            .I(N__36310));
    InMux I__6670 (
            .O(N__36313),
            .I(N__36307));
    LocalMux I__6669 (
            .O(N__36310),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ));
    LocalMux I__6668 (
            .O(N__36307),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ));
    InMux I__6667 (
            .O(N__36302),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ));
    InMux I__6666 (
            .O(N__36299),
            .I(N__36295));
    InMux I__6665 (
            .O(N__36298),
            .I(N__36292));
    LocalMux I__6664 (
            .O(N__36295),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ));
    LocalMux I__6663 (
            .O(N__36292),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ));
    InMux I__6662 (
            .O(N__36287),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ));
    InMux I__6661 (
            .O(N__36284),
            .I(N__36280));
    InMux I__6660 (
            .O(N__36283),
            .I(N__36277));
    LocalMux I__6659 (
            .O(N__36280),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ));
    LocalMux I__6658 (
            .O(N__36277),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ));
    InMux I__6657 (
            .O(N__36272),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ));
    InMux I__6656 (
            .O(N__36269),
            .I(N__36265));
    InMux I__6655 (
            .O(N__36268),
            .I(N__36262));
    LocalMux I__6654 (
            .O(N__36265),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ));
    LocalMux I__6653 (
            .O(N__36262),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ));
    InMux I__6652 (
            .O(N__36257),
            .I(bfn_13_10_0_));
    InMux I__6651 (
            .O(N__36254),
            .I(N__36250));
    InMux I__6650 (
            .O(N__36253),
            .I(N__36247));
    LocalMux I__6649 (
            .O(N__36250),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ));
    LocalMux I__6648 (
            .O(N__36247),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ));
    InMux I__6647 (
            .O(N__36242),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ));
    InMux I__6646 (
            .O(N__36239),
            .I(N__36235));
    InMux I__6645 (
            .O(N__36238),
            .I(N__36232));
    LocalMux I__6644 (
            .O(N__36235),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ));
    LocalMux I__6643 (
            .O(N__36232),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ));
    InMux I__6642 (
            .O(N__36227),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ));
    InMux I__6641 (
            .O(N__36224),
            .I(N__36220));
    InMux I__6640 (
            .O(N__36223),
            .I(N__36217));
    LocalMux I__6639 (
            .O(N__36220),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ));
    LocalMux I__6638 (
            .O(N__36217),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ));
    InMux I__6637 (
            .O(N__36212),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ));
    InMux I__6636 (
            .O(N__36209),
            .I(N__36205));
    InMux I__6635 (
            .O(N__36208),
            .I(N__36202));
    LocalMux I__6634 (
            .O(N__36205),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ));
    LocalMux I__6633 (
            .O(N__36202),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ));
    InMux I__6632 (
            .O(N__36197),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ));
    InMux I__6631 (
            .O(N__36194),
            .I(N__36190));
    InMux I__6630 (
            .O(N__36193),
            .I(N__36187));
    LocalMux I__6629 (
            .O(N__36190),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ));
    LocalMux I__6628 (
            .O(N__36187),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ));
    InMux I__6627 (
            .O(N__36182),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ));
    InMux I__6626 (
            .O(N__36179),
            .I(N__36175));
    InMux I__6625 (
            .O(N__36178),
            .I(N__36172));
    LocalMux I__6624 (
            .O(N__36175),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ));
    LocalMux I__6623 (
            .O(N__36172),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ));
    InMux I__6622 (
            .O(N__36167),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ));
    InMux I__6621 (
            .O(N__36164),
            .I(N__36161));
    LocalMux I__6620 (
            .O(N__36161),
            .I(N__36158));
    Odrv4 I__6619 (
            .O(N__36158),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ));
    InMux I__6618 (
            .O(N__36155),
            .I(N__36151));
    InMux I__6617 (
            .O(N__36154),
            .I(N__36148));
    LocalMux I__6616 (
            .O(N__36151),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ));
    LocalMux I__6615 (
            .O(N__36148),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ));
    InMux I__6614 (
            .O(N__36143),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ));
    InMux I__6613 (
            .O(N__36140),
            .I(N__36136));
    InMux I__6612 (
            .O(N__36139),
            .I(N__36133));
    LocalMux I__6611 (
            .O(N__36136),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ));
    LocalMux I__6610 (
            .O(N__36133),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ));
    InMux I__6609 (
            .O(N__36128),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ));
    InMux I__6608 (
            .O(N__36125),
            .I(N__36121));
    InMux I__6607 (
            .O(N__36124),
            .I(N__36118));
    LocalMux I__6606 (
            .O(N__36121),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ));
    LocalMux I__6605 (
            .O(N__36118),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ));
    InMux I__6604 (
            .O(N__36113),
            .I(bfn_13_9_0_));
    InMux I__6603 (
            .O(N__36110),
            .I(N__36106));
    InMux I__6602 (
            .O(N__36109),
            .I(N__36103));
    LocalMux I__6601 (
            .O(N__36106),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ));
    LocalMux I__6600 (
            .O(N__36103),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ));
    InMux I__6599 (
            .O(N__36098),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ));
    InMux I__6598 (
            .O(N__36095),
            .I(N__36092));
    LocalMux I__6597 (
            .O(N__36092),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ));
    InMux I__6596 (
            .O(N__36089),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ));
    InMux I__6595 (
            .O(N__36086),
            .I(N__36082));
    InMux I__6594 (
            .O(N__36085),
            .I(N__36079));
    LocalMux I__6593 (
            .O(N__36082),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ));
    LocalMux I__6592 (
            .O(N__36079),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ));
    InMux I__6591 (
            .O(N__36074),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ));
    InMux I__6590 (
            .O(N__36071),
            .I(N__36068));
    LocalMux I__6589 (
            .O(N__36068),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ));
    InMux I__6588 (
            .O(N__36065),
            .I(N__36061));
    InMux I__6587 (
            .O(N__36064),
            .I(N__36058));
    LocalMux I__6586 (
            .O(N__36061),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ));
    LocalMux I__6585 (
            .O(N__36058),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ));
    InMux I__6584 (
            .O(N__36053),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ));
    InMux I__6583 (
            .O(N__36050),
            .I(N__36046));
    InMux I__6582 (
            .O(N__36049),
            .I(N__36043));
    LocalMux I__6581 (
            .O(N__36046),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ));
    LocalMux I__6580 (
            .O(N__36043),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ));
    InMux I__6579 (
            .O(N__36038),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ));
    InMux I__6578 (
            .O(N__36035),
            .I(N__36031));
    InMux I__6577 (
            .O(N__36034),
            .I(N__36028));
    LocalMux I__6576 (
            .O(N__36031),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ));
    LocalMux I__6575 (
            .O(N__36028),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ));
    InMux I__6574 (
            .O(N__36023),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ));
    InMux I__6573 (
            .O(N__36020),
            .I(N__36016));
    InMux I__6572 (
            .O(N__36019),
            .I(N__36013));
    LocalMux I__6571 (
            .O(N__36016),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ));
    LocalMux I__6570 (
            .O(N__36013),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ));
    InMux I__6569 (
            .O(N__36008),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ));
    InMux I__6568 (
            .O(N__36005),
            .I(N__36001));
    InMux I__6567 (
            .O(N__36004),
            .I(N__35998));
    LocalMux I__6566 (
            .O(N__36001),
            .I(N__35993));
    LocalMux I__6565 (
            .O(N__35998),
            .I(N__35993));
    Odrv4 I__6564 (
            .O(N__35993),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ));
    InMux I__6563 (
            .O(N__35990),
            .I(bfn_13_8_0_));
    CascadeMux I__6562 (
            .O(N__35987),
            .I(N__35977));
    CascadeMux I__6561 (
            .O(N__35986),
            .I(N__35974));
    CascadeMux I__6560 (
            .O(N__35985),
            .I(N__35970));
    CascadeMux I__6559 (
            .O(N__35984),
            .I(N__35967));
    CascadeMux I__6558 (
            .O(N__35983),
            .I(N__35964));
    CascadeMux I__6557 (
            .O(N__35982),
            .I(N__35959));
    CascadeMux I__6556 (
            .O(N__35981),
            .I(N__35955));
    InMux I__6555 (
            .O(N__35980),
            .I(N__35952));
    InMux I__6554 (
            .O(N__35977),
            .I(N__35947));
    InMux I__6553 (
            .O(N__35974),
            .I(N__35947));
    InMux I__6552 (
            .O(N__35973),
            .I(N__35936));
    InMux I__6551 (
            .O(N__35970),
            .I(N__35936));
    InMux I__6550 (
            .O(N__35967),
            .I(N__35936));
    InMux I__6549 (
            .O(N__35964),
            .I(N__35936));
    InMux I__6548 (
            .O(N__35963),
            .I(N__35936));
    InMux I__6547 (
            .O(N__35962),
            .I(N__35927));
    InMux I__6546 (
            .O(N__35959),
            .I(N__35927));
    InMux I__6545 (
            .O(N__35958),
            .I(N__35927));
    InMux I__6544 (
            .O(N__35955),
            .I(N__35927));
    LocalMux I__6543 (
            .O(N__35952),
            .I(N__35924));
    LocalMux I__6542 (
            .O(N__35947),
            .I(N__35917));
    LocalMux I__6541 (
            .O(N__35936),
            .I(N__35917));
    LocalMux I__6540 (
            .O(N__35927),
            .I(N__35917));
    Span4Mux_v I__6539 (
            .O(N__35924),
            .I(N__35914));
    Span4Mux_v I__6538 (
            .O(N__35917),
            .I(N__35911));
    Sp12to4 I__6537 (
            .O(N__35914),
            .I(N__35906));
    Sp12to4 I__6536 (
            .O(N__35911),
            .I(N__35906));
    Span12Mux_h I__6535 (
            .O(N__35906),
            .I(N__35903));
    Odrv12 I__6534 (
            .O(N__35903),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    CascadeMux I__6533 (
            .O(N__35900),
            .I(N__35897));
    InMux I__6532 (
            .O(N__35897),
            .I(N__35894));
    LocalMux I__6531 (
            .O(N__35894),
            .I(N__35891));
    Span12Mux_v I__6530 (
            .O(N__35891),
            .I(N__35888));
    Span12Mux_h I__6529 (
            .O(N__35888),
            .I(N__35885));
    Odrv12 I__6528 (
            .O(N__35885),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    InMux I__6527 (
            .O(N__35882),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__6526 (
            .O(N__35879),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    IoInMux I__6525 (
            .O(N__35876),
            .I(N__35873));
    LocalMux I__6524 (
            .O(N__35873),
            .I(N__35870));
    Span4Mux_s0_v I__6523 (
            .O(N__35870),
            .I(N__35867));
    Odrv4 I__6522 (
            .O(N__35867),
            .I(GB_BUFFER_red_c_g_THRU_CO));
    InMux I__6521 (
            .O(N__35864),
            .I(N__35861));
    LocalMux I__6520 (
            .O(N__35861),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    CascadeMux I__6519 (
            .O(N__35858),
            .I(elapsed_time_ns_1_RNI24CN9_0_15_cascade_));
    InMux I__6518 (
            .O(N__35855),
            .I(N__35852));
    LocalMux I__6517 (
            .O(N__35852),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ));
    CascadeMux I__6516 (
            .O(N__35849),
            .I(N__35846));
    InMux I__6515 (
            .O(N__35846),
            .I(N__35843));
    LocalMux I__6514 (
            .O(N__35843),
            .I(N__35840));
    Sp12to4 I__6513 (
            .O(N__35840),
            .I(N__35837));
    Span12Mux_v I__6512 (
            .O(N__35837),
            .I(N__35834));
    Span12Mux_h I__6511 (
            .O(N__35834),
            .I(N__35831));
    Odrv12 I__6510 (
            .O(N__35831),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__6509 (
            .O(N__35828),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__6508 (
            .O(N__35825),
            .I(N__35822));
    LocalMux I__6507 (
            .O(N__35822),
            .I(N__35819));
    Span12Mux_v I__6506 (
            .O(N__35819),
            .I(N__35816));
    Span12Mux_h I__6505 (
            .O(N__35816),
            .I(N__35813));
    Odrv12 I__6504 (
            .O(N__35813),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__6503 (
            .O(N__35810),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    CascadeMux I__6502 (
            .O(N__35807),
            .I(N__35804));
    InMux I__6501 (
            .O(N__35804),
            .I(N__35801));
    LocalMux I__6500 (
            .O(N__35801),
            .I(N__35798));
    Span4Mux_v I__6499 (
            .O(N__35798),
            .I(N__35795));
    Sp12to4 I__6498 (
            .O(N__35795),
            .I(N__35792));
    Span12Mux_v I__6497 (
            .O(N__35792),
            .I(N__35789));
    Span12Mux_h I__6496 (
            .O(N__35789),
            .I(N__35786));
    Odrv12 I__6495 (
            .O(N__35786),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__6494 (
            .O(N__35783),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    CascadeMux I__6493 (
            .O(N__35780),
            .I(N__35777));
    InMux I__6492 (
            .O(N__35777),
            .I(N__35774));
    LocalMux I__6491 (
            .O(N__35774),
            .I(N__35771));
    Span12Mux_s11_v I__6490 (
            .O(N__35771),
            .I(N__35768));
    Span12Mux_h I__6489 (
            .O(N__35768),
            .I(N__35765));
    Odrv12 I__6488 (
            .O(N__35765),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__6487 (
            .O(N__35762),
            .I(bfn_12_24_0_));
    InMux I__6486 (
            .O(N__35759),
            .I(N__35756));
    LocalMux I__6485 (
            .O(N__35756),
            .I(N__35753));
    Span4Mux_v I__6484 (
            .O(N__35753),
            .I(N__35750));
    Sp12to4 I__6483 (
            .O(N__35750),
            .I(N__35747));
    Span12Mux_h I__6482 (
            .O(N__35747),
            .I(N__35744));
    Odrv12 I__6481 (
            .O(N__35744),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__6480 (
            .O(N__35741),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__6479 (
            .O(N__35738),
            .I(N__35735));
    LocalMux I__6478 (
            .O(N__35735),
            .I(N__35732));
    Span12Mux_v I__6477 (
            .O(N__35732),
            .I(N__35729));
    Span12Mux_h I__6476 (
            .O(N__35729),
            .I(N__35726));
    Odrv12 I__6475 (
            .O(N__35726),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__6474 (
            .O(N__35723),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__6473 (
            .O(N__35720),
            .I(N__35717));
    LocalMux I__6472 (
            .O(N__35717),
            .I(N__35714));
    Span12Mux_v I__6471 (
            .O(N__35714),
            .I(N__35711));
    Span12Mux_h I__6470 (
            .O(N__35711),
            .I(N__35708));
    Odrv12 I__6469 (
            .O(N__35708),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__6468 (
            .O(N__35705),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__6467 (
            .O(N__35702),
            .I(N__35699));
    LocalMux I__6466 (
            .O(N__35699),
            .I(N__35696));
    Span12Mux_v I__6465 (
            .O(N__35696),
            .I(N__35693));
    Span12Mux_h I__6464 (
            .O(N__35693),
            .I(N__35690));
    Odrv12 I__6463 (
            .O(N__35690),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__6462 (
            .O(N__35687),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__6461 (
            .O(N__35684),
            .I(N__35681));
    LocalMux I__6460 (
            .O(N__35681),
            .I(N__35678));
    Span12Mux_v I__6459 (
            .O(N__35678),
            .I(N__35675));
    Span12Mux_h I__6458 (
            .O(N__35675),
            .I(N__35672));
    Odrv12 I__6457 (
            .O(N__35672),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__6456 (
            .O(N__35669),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    CascadeMux I__6455 (
            .O(N__35666),
            .I(N__35663));
    InMux I__6454 (
            .O(N__35663),
            .I(N__35658));
    InMux I__6453 (
            .O(N__35662),
            .I(N__35655));
    InMux I__6452 (
            .O(N__35661),
            .I(N__35652));
    LocalMux I__6451 (
            .O(N__35658),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__6450 (
            .O(N__35655),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__6449 (
            .O(N__35652),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__6448 (
            .O(N__35645),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    CascadeMux I__6447 (
            .O(N__35642),
            .I(N__35638));
    InMux I__6446 (
            .O(N__35641),
            .I(N__35635));
    InMux I__6445 (
            .O(N__35638),
            .I(N__35632));
    LocalMux I__6444 (
            .O(N__35635),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__6443 (
            .O(N__35632),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__6442 (
            .O(N__35627),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__6441 (
            .O(N__35624),
            .I(N__35590));
    InMux I__6440 (
            .O(N__35623),
            .I(N__35590));
    InMux I__6439 (
            .O(N__35622),
            .I(N__35590));
    InMux I__6438 (
            .O(N__35621),
            .I(N__35590));
    InMux I__6437 (
            .O(N__35620),
            .I(N__35581));
    InMux I__6436 (
            .O(N__35619),
            .I(N__35581));
    InMux I__6435 (
            .O(N__35618),
            .I(N__35572));
    InMux I__6434 (
            .O(N__35617),
            .I(N__35572));
    InMux I__6433 (
            .O(N__35616),
            .I(N__35572));
    InMux I__6432 (
            .O(N__35615),
            .I(N__35572));
    InMux I__6431 (
            .O(N__35614),
            .I(N__35563));
    InMux I__6430 (
            .O(N__35613),
            .I(N__35563));
    InMux I__6429 (
            .O(N__35612),
            .I(N__35563));
    InMux I__6428 (
            .O(N__35611),
            .I(N__35563));
    InMux I__6427 (
            .O(N__35610),
            .I(N__35554));
    InMux I__6426 (
            .O(N__35609),
            .I(N__35554));
    InMux I__6425 (
            .O(N__35608),
            .I(N__35554));
    InMux I__6424 (
            .O(N__35607),
            .I(N__35554));
    InMux I__6423 (
            .O(N__35606),
            .I(N__35545));
    InMux I__6422 (
            .O(N__35605),
            .I(N__35545));
    InMux I__6421 (
            .O(N__35604),
            .I(N__35545));
    InMux I__6420 (
            .O(N__35603),
            .I(N__35545));
    InMux I__6419 (
            .O(N__35602),
            .I(N__35536));
    InMux I__6418 (
            .O(N__35601),
            .I(N__35536));
    InMux I__6417 (
            .O(N__35600),
            .I(N__35536));
    InMux I__6416 (
            .O(N__35599),
            .I(N__35536));
    LocalMux I__6415 (
            .O(N__35590),
            .I(N__35533));
    InMux I__6414 (
            .O(N__35589),
            .I(N__35524));
    InMux I__6413 (
            .O(N__35588),
            .I(N__35524));
    InMux I__6412 (
            .O(N__35587),
            .I(N__35524));
    InMux I__6411 (
            .O(N__35586),
            .I(N__35524));
    LocalMux I__6410 (
            .O(N__35581),
            .I(N__35519));
    LocalMux I__6409 (
            .O(N__35572),
            .I(N__35519));
    LocalMux I__6408 (
            .O(N__35563),
            .I(N__35510));
    LocalMux I__6407 (
            .O(N__35554),
            .I(N__35510));
    LocalMux I__6406 (
            .O(N__35545),
            .I(N__35510));
    LocalMux I__6405 (
            .O(N__35536),
            .I(N__35510));
    Span4Mux_h I__6404 (
            .O(N__35533),
            .I(N__35501));
    LocalMux I__6403 (
            .O(N__35524),
            .I(N__35501));
    Span4Mux_v I__6402 (
            .O(N__35519),
            .I(N__35501));
    Span4Mux_v I__6401 (
            .O(N__35510),
            .I(N__35501));
    Odrv4 I__6400 (
            .O(N__35501),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__6399 (
            .O(N__35498),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__6398 (
            .O(N__35495),
            .I(N__35491));
    InMux I__6397 (
            .O(N__35494),
            .I(N__35488));
    LocalMux I__6396 (
            .O(N__35491),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__6395 (
            .O(N__35488),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__6394 (
            .O(N__35483),
            .I(N__35479));
    CEMux I__6393 (
            .O(N__35482),
            .I(N__35476));
    LocalMux I__6392 (
            .O(N__35479),
            .I(N__35472));
    LocalMux I__6391 (
            .O(N__35476),
            .I(N__35469));
    CEMux I__6390 (
            .O(N__35475),
            .I(N__35466));
    Span4Mux_v I__6389 (
            .O(N__35472),
            .I(N__35459));
    Span4Mux_v I__6388 (
            .O(N__35469),
            .I(N__35459));
    LocalMux I__6387 (
            .O(N__35466),
            .I(N__35459));
    Span4Mux_v I__6386 (
            .O(N__35459),
            .I(N__35455));
    CEMux I__6385 (
            .O(N__35458),
            .I(N__35452));
    Span4Mux_v I__6384 (
            .O(N__35455),
            .I(N__35449));
    LocalMux I__6383 (
            .O(N__35452),
            .I(N__35446));
    Odrv4 I__6382 (
            .O(N__35449),
            .I(\delay_measurement_inst.delay_tr_timer.N_168_i ));
    Odrv12 I__6381 (
            .O(N__35446),
            .I(\delay_measurement_inst.delay_tr_timer.N_168_i ));
    InMux I__6380 (
            .O(N__35441),
            .I(N__35438));
    LocalMux I__6379 (
            .O(N__35438),
            .I(N__35435));
    Span4Mux_v I__6378 (
            .O(N__35435),
            .I(N__35432));
    Span4Mux_h I__6377 (
            .O(N__35432),
            .I(N__35429));
    Sp12to4 I__6376 (
            .O(N__35429),
            .I(N__35426));
    Span12Mux_v I__6375 (
            .O(N__35426),
            .I(N__35423));
    Odrv12 I__6374 (
            .O(N__35423),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__6373 (
            .O(N__35420),
            .I(N__35417));
    InMux I__6372 (
            .O(N__35417),
            .I(N__35414));
    LocalMux I__6371 (
            .O(N__35414),
            .I(N__35411));
    Span4Mux_v I__6370 (
            .O(N__35411),
            .I(N__35408));
    Span4Mux_h I__6369 (
            .O(N__35408),
            .I(N__35405));
    Sp12to4 I__6368 (
            .O(N__35405),
            .I(N__35402));
    Odrv12 I__6367 (
            .O(N__35402),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    InMux I__6366 (
            .O(N__35399),
            .I(N__35396));
    LocalMux I__6365 (
            .O(N__35396),
            .I(N__35393));
    Span4Mux_v I__6364 (
            .O(N__35393),
            .I(N__35390));
    Sp12to4 I__6363 (
            .O(N__35390),
            .I(N__35387));
    Span12Mux_h I__6362 (
            .O(N__35387),
            .I(N__35384));
    Odrv12 I__6361 (
            .O(N__35384),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    CascadeMux I__6360 (
            .O(N__35381),
            .I(N__35378));
    InMux I__6359 (
            .O(N__35378),
            .I(N__35375));
    LocalMux I__6358 (
            .O(N__35375),
            .I(N__35372));
    Span12Mux_v I__6357 (
            .O(N__35372),
            .I(N__35369));
    Span12Mux_h I__6356 (
            .O(N__35369),
            .I(N__35366));
    Odrv12 I__6355 (
            .O(N__35366),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    InMux I__6354 (
            .O(N__35363),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__6353 (
            .O(N__35360),
            .I(N__35357));
    LocalMux I__6352 (
            .O(N__35357),
            .I(N__35354));
    Span4Mux_v I__6351 (
            .O(N__35354),
            .I(N__35351));
    Sp12to4 I__6350 (
            .O(N__35351),
            .I(N__35348));
    Span12Mux_h I__6349 (
            .O(N__35348),
            .I(N__35345));
    Odrv12 I__6348 (
            .O(N__35345),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    CascadeMux I__6347 (
            .O(N__35342),
            .I(N__35339));
    InMux I__6346 (
            .O(N__35339),
            .I(N__35336));
    LocalMux I__6345 (
            .O(N__35336),
            .I(N__35333));
    Span12Mux_s10_v I__6344 (
            .O(N__35333),
            .I(N__35330));
    Span12Mux_h I__6343 (
            .O(N__35330),
            .I(N__35327));
    Odrv12 I__6342 (
            .O(N__35327),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    InMux I__6341 (
            .O(N__35324),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    InMux I__6340 (
            .O(N__35321),
            .I(N__35318));
    LocalMux I__6339 (
            .O(N__35318),
            .I(N__35315));
    Sp12to4 I__6338 (
            .O(N__35315),
            .I(N__35312));
    Span12Mux_s9_v I__6337 (
            .O(N__35312),
            .I(N__35309));
    Span12Mux_h I__6336 (
            .O(N__35309),
            .I(N__35306));
    Odrv12 I__6335 (
            .O(N__35306),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__6334 (
            .O(N__35303),
            .I(N__35300));
    InMux I__6333 (
            .O(N__35300),
            .I(N__35297));
    LocalMux I__6332 (
            .O(N__35297),
            .I(N__35294));
    Span4Mux_v I__6331 (
            .O(N__35294),
            .I(N__35291));
    Sp12to4 I__6330 (
            .O(N__35291),
            .I(N__35288));
    Span12Mux_h I__6329 (
            .O(N__35288),
            .I(N__35285));
    Odrv12 I__6328 (
            .O(N__35285),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__6327 (
            .O(N__35282),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    InMux I__6326 (
            .O(N__35279),
            .I(N__35276));
    LocalMux I__6325 (
            .O(N__35276),
            .I(N__35273));
    Span12Mux_s8_v I__6324 (
            .O(N__35273),
            .I(N__35270));
    Span12Mux_v I__6323 (
            .O(N__35270),
            .I(N__35267));
    Odrv12 I__6322 (
            .O(N__35267),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__6321 (
            .O(N__35264),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    CascadeMux I__6320 (
            .O(N__35261),
            .I(N__35258));
    InMux I__6319 (
            .O(N__35258),
            .I(N__35253));
    InMux I__6318 (
            .O(N__35257),
            .I(N__35250));
    InMux I__6317 (
            .O(N__35256),
            .I(N__35247));
    LocalMux I__6316 (
            .O(N__35253),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__6315 (
            .O(N__35250),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__6314 (
            .O(N__35247),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__6313 (
            .O(N__35240),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    CascadeMux I__6312 (
            .O(N__35237),
            .I(N__35234));
    InMux I__6311 (
            .O(N__35234),
            .I(N__35229));
    InMux I__6310 (
            .O(N__35233),
            .I(N__35226));
    InMux I__6309 (
            .O(N__35232),
            .I(N__35223));
    LocalMux I__6308 (
            .O(N__35229),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__6307 (
            .O(N__35226),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__6306 (
            .O(N__35223),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__6305 (
            .O(N__35216),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    CascadeMux I__6304 (
            .O(N__35213),
            .I(N__35210));
    InMux I__6303 (
            .O(N__35210),
            .I(N__35205));
    InMux I__6302 (
            .O(N__35209),
            .I(N__35202));
    InMux I__6301 (
            .O(N__35208),
            .I(N__35199));
    LocalMux I__6300 (
            .O(N__35205),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__6299 (
            .O(N__35202),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__6298 (
            .O(N__35199),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__6297 (
            .O(N__35192),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    CascadeMux I__6296 (
            .O(N__35189),
            .I(N__35186));
    InMux I__6295 (
            .O(N__35186),
            .I(N__35181));
    InMux I__6294 (
            .O(N__35185),
            .I(N__35178));
    InMux I__6293 (
            .O(N__35184),
            .I(N__35175));
    LocalMux I__6292 (
            .O(N__35181),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__6291 (
            .O(N__35178),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__6290 (
            .O(N__35175),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__6289 (
            .O(N__35168),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__6288 (
            .O(N__35165),
            .I(N__35162));
    InMux I__6287 (
            .O(N__35162),
            .I(N__35157));
    InMux I__6286 (
            .O(N__35161),
            .I(N__35154));
    InMux I__6285 (
            .O(N__35160),
            .I(N__35151));
    LocalMux I__6284 (
            .O(N__35157),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__6283 (
            .O(N__35154),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__6282 (
            .O(N__35151),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__6281 (
            .O(N__35144),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    CascadeMux I__6280 (
            .O(N__35141),
            .I(N__35138));
    InMux I__6279 (
            .O(N__35138),
            .I(N__35133));
    InMux I__6278 (
            .O(N__35137),
            .I(N__35130));
    InMux I__6277 (
            .O(N__35136),
            .I(N__35127));
    LocalMux I__6276 (
            .O(N__35133),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__6275 (
            .O(N__35130),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__6274 (
            .O(N__35127),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__6273 (
            .O(N__35120),
            .I(bfn_12_22_0_));
    CascadeMux I__6272 (
            .O(N__35117),
            .I(N__35114));
    InMux I__6271 (
            .O(N__35114),
            .I(N__35109));
    InMux I__6270 (
            .O(N__35113),
            .I(N__35106));
    InMux I__6269 (
            .O(N__35112),
            .I(N__35103));
    LocalMux I__6268 (
            .O(N__35109),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__6267 (
            .O(N__35106),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__6266 (
            .O(N__35103),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__6265 (
            .O(N__35096),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__6264 (
            .O(N__35093),
            .I(N__35088));
    InMux I__6263 (
            .O(N__35092),
            .I(N__35083));
    InMux I__6262 (
            .O(N__35091),
            .I(N__35083));
    LocalMux I__6261 (
            .O(N__35088),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__6260 (
            .O(N__35083),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__6259 (
            .O(N__35078),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    CascadeMux I__6258 (
            .O(N__35075),
            .I(N__35072));
    InMux I__6257 (
            .O(N__35072),
            .I(N__35067));
    InMux I__6256 (
            .O(N__35071),
            .I(N__35064));
    InMux I__6255 (
            .O(N__35070),
            .I(N__35061));
    LocalMux I__6254 (
            .O(N__35067),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__6253 (
            .O(N__35064),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__6252 (
            .O(N__35061),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__6251 (
            .O(N__35054),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    CascadeMux I__6250 (
            .O(N__35051),
            .I(N__35048));
    InMux I__6249 (
            .O(N__35048),
            .I(N__35043));
    InMux I__6248 (
            .O(N__35047),
            .I(N__35040));
    InMux I__6247 (
            .O(N__35046),
            .I(N__35037));
    LocalMux I__6246 (
            .O(N__35043),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__6245 (
            .O(N__35040),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__6244 (
            .O(N__35037),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__6243 (
            .O(N__35030),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    CascadeMux I__6242 (
            .O(N__35027),
            .I(N__35024));
    InMux I__6241 (
            .O(N__35024),
            .I(N__35019));
    InMux I__6240 (
            .O(N__35023),
            .I(N__35016));
    InMux I__6239 (
            .O(N__35022),
            .I(N__35013));
    LocalMux I__6238 (
            .O(N__35019),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__6237 (
            .O(N__35016),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__6236 (
            .O(N__35013),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__6235 (
            .O(N__35006),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    CascadeMux I__6234 (
            .O(N__35003),
            .I(N__35000));
    InMux I__6233 (
            .O(N__35000),
            .I(N__34995));
    InMux I__6232 (
            .O(N__34999),
            .I(N__34992));
    InMux I__6231 (
            .O(N__34998),
            .I(N__34989));
    LocalMux I__6230 (
            .O(N__34995),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__6229 (
            .O(N__34992),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__6228 (
            .O(N__34989),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__6227 (
            .O(N__34982),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__6226 (
            .O(N__34979),
            .I(N__34976));
    InMux I__6225 (
            .O(N__34976),
            .I(N__34971));
    InMux I__6224 (
            .O(N__34975),
            .I(N__34968));
    InMux I__6223 (
            .O(N__34974),
            .I(N__34965));
    LocalMux I__6222 (
            .O(N__34971),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__6221 (
            .O(N__34968),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__6220 (
            .O(N__34965),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__6219 (
            .O(N__34958),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    CascadeMux I__6218 (
            .O(N__34955),
            .I(N__34952));
    InMux I__6217 (
            .O(N__34952),
            .I(N__34947));
    InMux I__6216 (
            .O(N__34951),
            .I(N__34944));
    InMux I__6215 (
            .O(N__34950),
            .I(N__34941));
    LocalMux I__6214 (
            .O(N__34947),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__6213 (
            .O(N__34944),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__6212 (
            .O(N__34941),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__6211 (
            .O(N__34934),
            .I(bfn_12_21_0_));
    CascadeMux I__6210 (
            .O(N__34931),
            .I(N__34928));
    InMux I__6209 (
            .O(N__34928),
            .I(N__34923));
    InMux I__6208 (
            .O(N__34927),
            .I(N__34920));
    InMux I__6207 (
            .O(N__34926),
            .I(N__34917));
    LocalMux I__6206 (
            .O(N__34923),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__6205 (
            .O(N__34920),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__6204 (
            .O(N__34917),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__6203 (
            .O(N__34910),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__6202 (
            .O(N__34907),
            .I(N__34904));
    InMux I__6201 (
            .O(N__34904),
            .I(N__34899));
    InMux I__6200 (
            .O(N__34903),
            .I(N__34896));
    InMux I__6199 (
            .O(N__34902),
            .I(N__34893));
    LocalMux I__6198 (
            .O(N__34899),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__6197 (
            .O(N__34896),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__6196 (
            .O(N__34893),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__6195 (
            .O(N__34886),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__6194 (
            .O(N__34883),
            .I(N__34878));
    InMux I__6193 (
            .O(N__34882),
            .I(N__34873));
    InMux I__6192 (
            .O(N__34881),
            .I(N__34873));
    LocalMux I__6191 (
            .O(N__34878),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__6190 (
            .O(N__34873),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__6189 (
            .O(N__34868),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    CascadeMux I__6188 (
            .O(N__34865),
            .I(N__34862));
    InMux I__6187 (
            .O(N__34862),
            .I(N__34857));
    InMux I__6186 (
            .O(N__34861),
            .I(N__34854));
    InMux I__6185 (
            .O(N__34860),
            .I(N__34851));
    LocalMux I__6184 (
            .O(N__34857),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__6183 (
            .O(N__34854),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__6182 (
            .O(N__34851),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__6181 (
            .O(N__34844),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    CascadeMux I__6180 (
            .O(N__34841),
            .I(N__34836));
    CascadeMux I__6179 (
            .O(N__34840),
            .I(N__34833));
    InMux I__6178 (
            .O(N__34839),
            .I(N__34830));
    InMux I__6177 (
            .O(N__34836),
            .I(N__34825));
    InMux I__6176 (
            .O(N__34833),
            .I(N__34825));
    LocalMux I__6175 (
            .O(N__34830),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__6174 (
            .O(N__34825),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__6173 (
            .O(N__34820),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__6172 (
            .O(N__34817),
            .I(N__34814));
    InMux I__6171 (
            .O(N__34814),
            .I(N__34809));
    InMux I__6170 (
            .O(N__34813),
            .I(N__34806));
    InMux I__6169 (
            .O(N__34812),
            .I(N__34803));
    LocalMux I__6168 (
            .O(N__34809),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__6167 (
            .O(N__34806),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__6166 (
            .O(N__34803),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__6165 (
            .O(N__34796),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__6164 (
            .O(N__34793),
            .I(N__34790));
    InMux I__6163 (
            .O(N__34790),
            .I(N__34785));
    InMux I__6162 (
            .O(N__34789),
            .I(N__34782));
    InMux I__6161 (
            .O(N__34788),
            .I(N__34779));
    LocalMux I__6160 (
            .O(N__34785),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__6159 (
            .O(N__34782),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__6158 (
            .O(N__34779),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__6157 (
            .O(N__34772),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__6156 (
            .O(N__34769),
            .I(N__34766));
    InMux I__6155 (
            .O(N__34766),
            .I(N__34761));
    InMux I__6154 (
            .O(N__34765),
            .I(N__34758));
    InMux I__6153 (
            .O(N__34764),
            .I(N__34755));
    LocalMux I__6152 (
            .O(N__34761),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__6151 (
            .O(N__34758),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__6150 (
            .O(N__34755),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__6149 (
            .O(N__34748),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    CascadeMux I__6148 (
            .O(N__34745),
            .I(N__34742));
    InMux I__6147 (
            .O(N__34742),
            .I(N__34737));
    InMux I__6146 (
            .O(N__34741),
            .I(N__34734));
    InMux I__6145 (
            .O(N__34740),
            .I(N__34731));
    LocalMux I__6144 (
            .O(N__34737),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__6143 (
            .O(N__34734),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__6142 (
            .O(N__34731),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__6141 (
            .O(N__34724),
            .I(bfn_12_20_0_));
    CascadeMux I__6140 (
            .O(N__34721),
            .I(N__34718));
    InMux I__6139 (
            .O(N__34718),
            .I(N__34713));
    InMux I__6138 (
            .O(N__34717),
            .I(N__34710));
    InMux I__6137 (
            .O(N__34716),
            .I(N__34707));
    LocalMux I__6136 (
            .O(N__34713),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__6135 (
            .O(N__34710),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__6134 (
            .O(N__34707),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__6133 (
            .O(N__34700),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__6132 (
            .O(N__34697),
            .I(N__34694));
    InMux I__6131 (
            .O(N__34694),
            .I(N__34689));
    InMux I__6130 (
            .O(N__34693),
            .I(N__34686));
    InMux I__6129 (
            .O(N__34692),
            .I(N__34683));
    LocalMux I__6128 (
            .O(N__34689),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__6127 (
            .O(N__34686),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__6126 (
            .O(N__34683),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__6125 (
            .O(N__34676),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__6124 (
            .O(N__34673),
            .I(N__34670));
    LocalMux I__6123 (
            .O(N__34670),
            .I(N__34666));
    InMux I__6122 (
            .O(N__34669),
            .I(N__34663));
    Odrv12 I__6121 (
            .O(N__34666),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_17));
    LocalMux I__6120 (
            .O(N__34663),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_17));
    InMux I__6119 (
            .O(N__34658),
            .I(N__34652));
    InMux I__6118 (
            .O(N__34657),
            .I(N__34652));
    LocalMux I__6117 (
            .O(N__34652),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ));
    InMux I__6116 (
            .O(N__34649),
            .I(N__34646));
    LocalMux I__6115 (
            .O(N__34646),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt18 ));
    InMux I__6114 (
            .O(N__34643),
            .I(N__34639));
    InMux I__6113 (
            .O(N__34642),
            .I(N__34636));
    LocalMux I__6112 (
            .O(N__34639),
            .I(N__34633));
    LocalMux I__6111 (
            .O(N__34636),
            .I(N__34630));
    Odrv12 I__6110 (
            .O(N__34633),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_18));
    Odrv4 I__6109 (
            .O(N__34630),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_18));
    InMux I__6108 (
            .O(N__34625),
            .I(N__34619));
    InMux I__6107 (
            .O(N__34624),
            .I(N__34619));
    LocalMux I__6106 (
            .O(N__34619),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ));
    InMux I__6105 (
            .O(N__34616),
            .I(N__34610));
    InMux I__6104 (
            .O(N__34615),
            .I(N__34610));
    LocalMux I__6103 (
            .O(N__34610),
            .I(N__34607));
    Odrv4 I__6102 (
            .O(N__34607),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ));
    CascadeMux I__6101 (
            .O(N__34604),
            .I(N__34600));
    CascadeMux I__6100 (
            .O(N__34603),
            .I(N__34597));
    InMux I__6099 (
            .O(N__34600),
            .I(N__34592));
    InMux I__6098 (
            .O(N__34597),
            .I(N__34592));
    LocalMux I__6097 (
            .O(N__34592),
            .I(N__34588));
    InMux I__6096 (
            .O(N__34591),
            .I(N__34585));
    Span4Mux_h I__6095 (
            .O(N__34588),
            .I(N__34582));
    LocalMux I__6094 (
            .O(N__34585),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ));
    Odrv4 I__6093 (
            .O(N__34582),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ));
    InMux I__6092 (
            .O(N__34577),
            .I(N__34571));
    InMux I__6091 (
            .O(N__34576),
            .I(N__34571));
    LocalMux I__6090 (
            .O(N__34571),
            .I(N__34567));
    InMux I__6089 (
            .O(N__34570),
            .I(N__34564));
    Span4Mux_h I__6088 (
            .O(N__34567),
            .I(N__34561));
    LocalMux I__6087 (
            .O(N__34564),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ));
    Odrv4 I__6086 (
            .O(N__34561),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ));
    CascadeMux I__6085 (
            .O(N__34556),
            .I(N__34553));
    InMux I__6084 (
            .O(N__34553),
            .I(N__34550));
    LocalMux I__6083 (
            .O(N__34550),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ));
    CascadeMux I__6082 (
            .O(N__34547),
            .I(N__34540));
    InMux I__6081 (
            .O(N__34546),
            .I(N__34537));
    InMux I__6080 (
            .O(N__34545),
            .I(N__34534));
    InMux I__6079 (
            .O(N__34544),
            .I(N__34531));
    InMux I__6078 (
            .O(N__34543),
            .I(N__34528));
    InMux I__6077 (
            .O(N__34540),
            .I(N__34524));
    LocalMux I__6076 (
            .O(N__34537),
            .I(N__34517));
    LocalMux I__6075 (
            .O(N__34534),
            .I(N__34517));
    LocalMux I__6074 (
            .O(N__34531),
            .I(N__34517));
    LocalMux I__6073 (
            .O(N__34528),
            .I(N__34514));
    InMux I__6072 (
            .O(N__34527),
            .I(N__34511));
    LocalMux I__6071 (
            .O(N__34524),
            .I(N__34506));
    Span4Mux_v I__6070 (
            .O(N__34517),
            .I(N__34506));
    Span4Mux_v I__6069 (
            .O(N__34514),
            .I(N__34503));
    LocalMux I__6068 (
            .O(N__34511),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__6067 (
            .O(N__34506),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__6066 (
            .O(N__34503),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__6065 (
            .O(N__34496),
            .I(N__34472));
    InMux I__6064 (
            .O(N__34495),
            .I(N__34472));
    InMux I__6063 (
            .O(N__34494),
            .I(N__34472));
    InMux I__6062 (
            .O(N__34493),
            .I(N__34472));
    InMux I__6061 (
            .O(N__34492),
            .I(N__34463));
    InMux I__6060 (
            .O(N__34491),
            .I(N__34463));
    InMux I__6059 (
            .O(N__34490),
            .I(N__34463));
    InMux I__6058 (
            .O(N__34489),
            .I(N__34463));
    InMux I__6057 (
            .O(N__34488),
            .I(N__34446));
    InMux I__6056 (
            .O(N__34487),
            .I(N__34446));
    InMux I__6055 (
            .O(N__34486),
            .I(N__34446));
    InMux I__6054 (
            .O(N__34485),
            .I(N__34446));
    InMux I__6053 (
            .O(N__34484),
            .I(N__34437));
    InMux I__6052 (
            .O(N__34483),
            .I(N__34437));
    InMux I__6051 (
            .O(N__34482),
            .I(N__34437));
    InMux I__6050 (
            .O(N__34481),
            .I(N__34437));
    LocalMux I__6049 (
            .O(N__34472),
            .I(N__34428));
    LocalMux I__6048 (
            .O(N__34463),
            .I(N__34428));
    InMux I__6047 (
            .O(N__34462),
            .I(N__34421));
    InMux I__6046 (
            .O(N__34461),
            .I(N__34421));
    InMux I__6045 (
            .O(N__34460),
            .I(N__34421));
    InMux I__6044 (
            .O(N__34459),
            .I(N__34410));
    InMux I__6043 (
            .O(N__34458),
            .I(N__34410));
    InMux I__6042 (
            .O(N__34457),
            .I(N__34410));
    InMux I__6041 (
            .O(N__34456),
            .I(N__34410));
    InMux I__6040 (
            .O(N__34455),
            .I(N__34410));
    LocalMux I__6039 (
            .O(N__34446),
            .I(N__34401));
    LocalMux I__6038 (
            .O(N__34437),
            .I(N__34401));
    InMux I__6037 (
            .O(N__34436),
            .I(N__34392));
    InMux I__6036 (
            .O(N__34435),
            .I(N__34392));
    InMux I__6035 (
            .O(N__34434),
            .I(N__34392));
    InMux I__6034 (
            .O(N__34433),
            .I(N__34392));
    Span4Mux_v I__6033 (
            .O(N__34428),
            .I(N__34387));
    LocalMux I__6032 (
            .O(N__34421),
            .I(N__34387));
    LocalMux I__6031 (
            .O(N__34410),
            .I(N__34384));
    InMux I__6030 (
            .O(N__34409),
            .I(N__34375));
    InMux I__6029 (
            .O(N__34408),
            .I(N__34375));
    InMux I__6028 (
            .O(N__34407),
            .I(N__34375));
    InMux I__6027 (
            .O(N__34406),
            .I(N__34375));
    Span4Mux_h I__6026 (
            .O(N__34401),
            .I(N__34366));
    LocalMux I__6025 (
            .O(N__34392),
            .I(N__34366));
    Span4Mux_v I__6024 (
            .O(N__34387),
            .I(N__34366));
    Span4Mux_v I__6023 (
            .O(N__34384),
            .I(N__34366));
    LocalMux I__6022 (
            .O(N__34375),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    Odrv4 I__6021 (
            .O(N__34366),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    InMux I__6020 (
            .O(N__34361),
            .I(N__34355));
    InMux I__6019 (
            .O(N__34360),
            .I(N__34348));
    InMux I__6018 (
            .O(N__34359),
            .I(N__34348));
    InMux I__6017 (
            .O(N__34358),
            .I(N__34348));
    LocalMux I__6016 (
            .O(N__34355),
            .I(N__34345));
    LocalMux I__6015 (
            .O(N__34348),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__6014 (
            .O(N__34345),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__6013 (
            .O(N__34340),
            .I(N__34337));
    LocalMux I__6012 (
            .O(N__34337),
            .I(N__34334));
    Span4Mux_h I__6011 (
            .O(N__34334),
            .I(N__34330));
    CascadeMux I__6010 (
            .O(N__34333),
            .I(N__34327));
    Span4Mux_v I__6009 (
            .O(N__34330),
            .I(N__34323));
    InMux I__6008 (
            .O(N__34327),
            .I(N__34320));
    InMux I__6007 (
            .O(N__34326),
            .I(N__34317));
    Odrv4 I__6006 (
            .O(N__34323),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__6005 (
            .O(N__34320),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__6004 (
            .O(N__34317),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__6003 (
            .O(N__34310),
            .I(bfn_12_19_0_));
    InMux I__6002 (
            .O(N__34307),
            .I(N__34304));
    LocalMux I__6001 (
            .O(N__34304),
            .I(N__34301));
    Span4Mux_v I__6000 (
            .O(N__34301),
            .I(N__34298));
    Span4Mux_v I__5999 (
            .O(N__34298),
            .I(N__34294));
    CascadeMux I__5998 (
            .O(N__34297),
            .I(N__34291));
    Span4Mux_h I__5997 (
            .O(N__34294),
            .I(N__34287));
    InMux I__5996 (
            .O(N__34291),
            .I(N__34284));
    InMux I__5995 (
            .O(N__34290),
            .I(N__34281));
    Odrv4 I__5994 (
            .O(N__34287),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__5993 (
            .O(N__34284),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__5992 (
            .O(N__34281),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__5991 (
            .O(N__34274),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CEMux I__5990 (
            .O(N__34271),
            .I(N__34266));
    CEMux I__5989 (
            .O(N__34270),
            .I(N__34263));
    CEMux I__5988 (
            .O(N__34269),
            .I(N__34260));
    LocalMux I__5987 (
            .O(N__34266),
            .I(N__34256));
    LocalMux I__5986 (
            .O(N__34263),
            .I(N__34251));
    LocalMux I__5985 (
            .O(N__34260),
            .I(N__34251));
    CEMux I__5984 (
            .O(N__34259),
            .I(N__34248));
    Span4Mux_v I__5983 (
            .O(N__34256),
            .I(N__34241));
    Span4Mux_v I__5982 (
            .O(N__34251),
            .I(N__34241));
    LocalMux I__5981 (
            .O(N__34248),
            .I(N__34238));
    CEMux I__5980 (
            .O(N__34247),
            .I(N__34235));
    CEMux I__5979 (
            .O(N__34246),
            .I(N__34232));
    Span4Mux_v I__5978 (
            .O(N__34241),
            .I(N__34227));
    Span4Mux_v I__5977 (
            .O(N__34238),
            .I(N__34227));
    LocalMux I__5976 (
            .O(N__34235),
            .I(N__34224));
    LocalMux I__5975 (
            .O(N__34232),
            .I(N__34221));
    Span4Mux_v I__5974 (
            .O(N__34227),
            .I(N__34218));
    Span4Mux_v I__5973 (
            .O(N__34224),
            .I(N__34215));
    Span4Mux_h I__5972 (
            .O(N__34221),
            .I(N__34212));
    Odrv4 I__5971 (
            .O(N__34218),
            .I(\delay_measurement_inst.delay_tr_timer.N_167_i ));
    Odrv4 I__5970 (
            .O(N__34215),
            .I(\delay_measurement_inst.delay_tr_timer.N_167_i ));
    Odrv4 I__5969 (
            .O(N__34212),
            .I(\delay_measurement_inst.delay_tr_timer.N_167_i ));
    InMux I__5968 (
            .O(N__34205),
            .I(N__34202));
    LocalMux I__5967 (
            .O(N__34202),
            .I(N__34199));
    Span4Mux_h I__5966 (
            .O(N__34199),
            .I(N__34194));
    InMux I__5965 (
            .O(N__34198),
            .I(N__34191));
    InMux I__5964 (
            .O(N__34197),
            .I(N__34188));
    Odrv4 I__5963 (
            .O(N__34194),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__5962 (
            .O(N__34191),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__5961 (
            .O(N__34188),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    CascadeMux I__5960 (
            .O(N__34181),
            .I(\phase_controller_inst1.stoper_hc.un4_start_0_cascade_ ));
    InMux I__5959 (
            .O(N__34178),
            .I(N__34175));
    LocalMux I__5958 (
            .O(N__34175),
            .I(N__34171));
    InMux I__5957 (
            .O(N__34174),
            .I(N__34168));
    Span4Mux_h I__5956 (
            .O(N__34171),
            .I(N__34162));
    LocalMux I__5955 (
            .O(N__34168),
            .I(N__34162));
    InMux I__5954 (
            .O(N__34167),
            .I(N__34159));
    Odrv4 I__5953 (
            .O(N__34162),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ));
    LocalMux I__5952 (
            .O(N__34159),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ));
    CascadeMux I__5951 (
            .O(N__34154),
            .I(N__34150));
    InMux I__5950 (
            .O(N__34153),
            .I(N__34145));
    InMux I__5949 (
            .O(N__34150),
            .I(N__34145));
    LocalMux I__5948 (
            .O(N__34145),
            .I(N__34140));
    InMux I__5947 (
            .O(N__34144),
            .I(N__34137));
    InMux I__5946 (
            .O(N__34143),
            .I(N__34134));
    Span4Mux_v I__5945 (
            .O(N__34140),
            .I(N__34129));
    LocalMux I__5944 (
            .O(N__34137),
            .I(N__34129));
    LocalMux I__5943 (
            .O(N__34134),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__5942 (
            .O(N__34129),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__5941 (
            .O(N__34124),
            .I(N__34120));
    InMux I__5940 (
            .O(N__34123),
            .I(N__34117));
    LocalMux I__5939 (
            .O(N__34120),
            .I(N__34113));
    LocalMux I__5938 (
            .O(N__34117),
            .I(N__34110));
    InMux I__5937 (
            .O(N__34116),
            .I(N__34107));
    Span4Mux_v I__5936 (
            .O(N__34113),
            .I(N__34102));
    Span4Mux_h I__5935 (
            .O(N__34110),
            .I(N__34102));
    LocalMux I__5934 (
            .O(N__34107),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ));
    Odrv4 I__5933 (
            .O(N__34102),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ));
    InMux I__5932 (
            .O(N__34097),
            .I(N__34094));
    LocalMux I__5931 (
            .O(N__34094),
            .I(N__34090));
    InMux I__5930 (
            .O(N__34093),
            .I(N__34087));
    Span4Mux_v I__5929 (
            .O(N__34090),
            .I(N__34081));
    LocalMux I__5928 (
            .O(N__34087),
            .I(N__34081));
    InMux I__5927 (
            .O(N__34086),
            .I(N__34078));
    Span4Mux_h I__5926 (
            .O(N__34081),
            .I(N__34075));
    LocalMux I__5925 (
            .O(N__34078),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ));
    Odrv4 I__5924 (
            .O(N__34075),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ));
    InMux I__5923 (
            .O(N__34070),
            .I(N__34067));
    LocalMux I__5922 (
            .O(N__34067),
            .I(N__34064));
    Span4Mux_v I__5921 (
            .O(N__34064),
            .I(N__34058));
    InMux I__5920 (
            .O(N__34063),
            .I(N__34051));
    InMux I__5919 (
            .O(N__34062),
            .I(N__34051));
    InMux I__5918 (
            .O(N__34061),
            .I(N__34051));
    Span4Mux_h I__5917 (
            .O(N__34058),
            .I(N__34046));
    LocalMux I__5916 (
            .O(N__34051),
            .I(N__34046));
    Odrv4 I__5915 (
            .O(N__34046),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ));
    InMux I__5914 (
            .O(N__34043),
            .I(N__34040));
    LocalMux I__5913 (
            .O(N__34040),
            .I(N__34037));
    Span4Mux_h I__5912 (
            .O(N__34037),
            .I(N__34034));
    Odrv4 I__5911 (
            .O(N__34034),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ));
    InMux I__5910 (
            .O(N__34031),
            .I(N__34027));
    InMux I__5909 (
            .O(N__34030),
            .I(N__34024));
    LocalMux I__5908 (
            .O(N__34027),
            .I(N__34018));
    LocalMux I__5907 (
            .O(N__34024),
            .I(N__34014));
    InMux I__5906 (
            .O(N__34023),
            .I(N__34007));
    InMux I__5905 (
            .O(N__34022),
            .I(N__34007));
    InMux I__5904 (
            .O(N__34021),
            .I(N__34007));
    Span4Mux_v I__5903 (
            .O(N__34018),
            .I(N__34004));
    InMux I__5902 (
            .O(N__34017),
            .I(N__34001));
    Span4Mux_h I__5901 (
            .O(N__34014),
            .I(N__33998));
    LocalMux I__5900 (
            .O(N__34007),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__5899 (
            .O(N__34004),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__5898 (
            .O(N__34001),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__5897 (
            .O(N__33998),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__5896 (
            .O(N__33989),
            .I(N__33986));
    LocalMux I__5895 (
            .O(N__33986),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt16 ));
    InMux I__5894 (
            .O(N__33983),
            .I(N__33979));
    InMux I__5893 (
            .O(N__33982),
            .I(N__33976));
    LocalMux I__5892 (
            .O(N__33979),
            .I(N__33973));
    LocalMux I__5891 (
            .O(N__33976),
            .I(N__33970));
    Odrv12 I__5890 (
            .O(N__33973),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_16));
    Odrv4 I__5889 (
            .O(N__33970),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_16));
    InMux I__5888 (
            .O(N__33965),
            .I(N__33959));
    InMux I__5887 (
            .O(N__33964),
            .I(N__33959));
    LocalMux I__5886 (
            .O(N__33959),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ));
    InMux I__5885 (
            .O(N__33956),
            .I(N__33950));
    InMux I__5884 (
            .O(N__33955),
            .I(N__33950));
    LocalMux I__5883 (
            .O(N__33950),
            .I(N__33946));
    InMux I__5882 (
            .O(N__33949),
            .I(N__33943));
    Span4Mux_h I__5881 (
            .O(N__33946),
            .I(N__33940));
    LocalMux I__5880 (
            .O(N__33943),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ));
    Odrv4 I__5879 (
            .O(N__33940),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ));
    CascadeMux I__5878 (
            .O(N__33935),
            .I(N__33931));
    CascadeMux I__5877 (
            .O(N__33934),
            .I(N__33928));
    InMux I__5876 (
            .O(N__33931),
            .I(N__33923));
    InMux I__5875 (
            .O(N__33928),
            .I(N__33923));
    LocalMux I__5874 (
            .O(N__33923),
            .I(N__33919));
    InMux I__5873 (
            .O(N__33922),
            .I(N__33916));
    Span4Mux_h I__5872 (
            .O(N__33919),
            .I(N__33913));
    LocalMux I__5871 (
            .O(N__33916),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ));
    Odrv4 I__5870 (
            .O(N__33913),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ));
    CascadeMux I__5869 (
            .O(N__33908),
            .I(N__33905));
    InMux I__5868 (
            .O(N__33905),
            .I(N__33902));
    LocalMux I__5867 (
            .O(N__33902),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ));
    InMux I__5866 (
            .O(N__33899),
            .I(N__33896));
    LocalMux I__5865 (
            .O(N__33896),
            .I(N__33892));
    InMux I__5864 (
            .O(N__33895),
            .I(N__33889));
    Span4Mux_v I__5863 (
            .O(N__33892),
            .I(N__33884));
    LocalMux I__5862 (
            .O(N__33889),
            .I(N__33884));
    Odrv4 I__5861 (
            .O(N__33884),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_2));
    InMux I__5860 (
            .O(N__33881),
            .I(N__33878));
    LocalMux I__5859 (
            .O(N__33878),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ));
    InMux I__5858 (
            .O(N__33875),
            .I(N__33871));
    InMux I__5857 (
            .O(N__33874),
            .I(N__33868));
    LocalMux I__5856 (
            .O(N__33871),
            .I(N__33865));
    LocalMux I__5855 (
            .O(N__33868),
            .I(N__33862));
    Odrv12 I__5854 (
            .O(N__33865),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_6));
    Odrv4 I__5853 (
            .O(N__33862),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_6));
    CascadeMux I__5852 (
            .O(N__33857),
            .I(N__33854));
    InMux I__5851 (
            .O(N__33854),
            .I(N__33851));
    LocalMux I__5850 (
            .O(N__33851),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ));
    InMux I__5849 (
            .O(N__33848),
            .I(N__33845));
    LocalMux I__5848 (
            .O(N__33845),
            .I(N__33841));
    InMux I__5847 (
            .O(N__33844),
            .I(N__33838));
    Odrv4 I__5846 (
            .O(N__33841),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_19));
    LocalMux I__5845 (
            .O(N__33838),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_19));
    InMux I__5844 (
            .O(N__33833),
            .I(N__33830));
    LocalMux I__5843 (
            .O(N__33830),
            .I(N__33826));
    InMux I__5842 (
            .O(N__33829),
            .I(N__33823));
    Span4Mux_v I__5841 (
            .O(N__33826),
            .I(N__33818));
    LocalMux I__5840 (
            .O(N__33823),
            .I(N__33818));
    Odrv4 I__5839 (
            .O(N__33818),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_3));
    InMux I__5838 (
            .O(N__33815),
            .I(N__33812));
    LocalMux I__5837 (
            .O(N__33812),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ));
    InMux I__5836 (
            .O(N__33809),
            .I(N__33805));
    InMux I__5835 (
            .O(N__33808),
            .I(N__33802));
    LocalMux I__5834 (
            .O(N__33805),
            .I(N__33799));
    LocalMux I__5833 (
            .O(N__33802),
            .I(N__33796));
    Odrv12 I__5832 (
            .O(N__33799),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_7));
    Odrv4 I__5831 (
            .O(N__33796),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_7));
    CascadeMux I__5830 (
            .O(N__33791),
            .I(N__33788));
    InMux I__5829 (
            .O(N__33788),
            .I(N__33785));
    LocalMux I__5828 (
            .O(N__33785),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ));
    InMux I__5827 (
            .O(N__33782),
            .I(N__33778));
    InMux I__5826 (
            .O(N__33781),
            .I(N__33775));
    LocalMux I__5825 (
            .O(N__33778),
            .I(N__33772));
    LocalMux I__5824 (
            .O(N__33775),
            .I(N__33769));
    Odrv4 I__5823 (
            .O(N__33772),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_10));
    Odrv4 I__5822 (
            .O(N__33769),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_10));
    InMux I__5821 (
            .O(N__33764),
            .I(N__33761));
    LocalMux I__5820 (
            .O(N__33761),
            .I(N__33758));
    Odrv4 I__5819 (
            .O(N__33758),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ));
    InMux I__5818 (
            .O(N__33755),
            .I(N__33751));
    InMux I__5817 (
            .O(N__33754),
            .I(N__33748));
    LocalMux I__5816 (
            .O(N__33751),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_25));
    LocalMux I__5815 (
            .O(N__33748),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_25));
    InMux I__5814 (
            .O(N__33743),
            .I(N__33737));
    InMux I__5813 (
            .O(N__33742),
            .I(N__33737));
    LocalMux I__5812 (
            .O(N__33737),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ));
    InMux I__5811 (
            .O(N__33734),
            .I(N__33730));
    InMux I__5810 (
            .O(N__33733),
            .I(N__33727));
    LocalMux I__5809 (
            .O(N__33730),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_22));
    LocalMux I__5808 (
            .O(N__33727),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_22));
    InMux I__5807 (
            .O(N__33722),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ));
    InMux I__5806 (
            .O(N__33719),
            .I(N__33715));
    InMux I__5805 (
            .O(N__33718),
            .I(N__33712));
    LocalMux I__5804 (
            .O(N__33715),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_23));
    LocalMux I__5803 (
            .O(N__33712),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_23));
    InMux I__5802 (
            .O(N__33707),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ));
    InMux I__5801 (
            .O(N__33704),
            .I(N__33700));
    InMux I__5800 (
            .O(N__33703),
            .I(N__33697));
    LocalMux I__5799 (
            .O(N__33700),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_24));
    LocalMux I__5798 (
            .O(N__33697),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_24));
    InMux I__5797 (
            .O(N__33692),
            .I(bfn_12_10_0_));
    InMux I__5796 (
            .O(N__33689),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ));
    InMux I__5795 (
            .O(N__33686),
            .I(N__33682));
    InMux I__5794 (
            .O(N__33685),
            .I(N__33679));
    LocalMux I__5793 (
            .O(N__33682),
            .I(N__33676));
    LocalMux I__5792 (
            .O(N__33679),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_26));
    Odrv4 I__5791 (
            .O(N__33676),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_26));
    InMux I__5790 (
            .O(N__33671),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ));
    InMux I__5789 (
            .O(N__33668),
            .I(N__33664));
    InMux I__5788 (
            .O(N__33667),
            .I(N__33661));
    LocalMux I__5787 (
            .O(N__33664),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_27));
    LocalMux I__5786 (
            .O(N__33661),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_27));
    InMux I__5785 (
            .O(N__33656),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ));
    InMux I__5784 (
            .O(N__33653),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ));
    InMux I__5783 (
            .O(N__33650),
            .I(N__33646));
    InMux I__5782 (
            .O(N__33649),
            .I(N__33643));
    LocalMux I__5781 (
            .O(N__33646),
            .I(N__33640));
    LocalMux I__5780 (
            .O(N__33643),
            .I(N__33637));
    Odrv12 I__5779 (
            .O(N__33640),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_4));
    Odrv4 I__5778 (
            .O(N__33637),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_4));
    InMux I__5777 (
            .O(N__33632),
            .I(N__33629));
    LocalMux I__5776 (
            .O(N__33629),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ));
    InMux I__5775 (
            .O(N__33626),
            .I(N__33623));
    LocalMux I__5774 (
            .O(N__33623),
            .I(N__33619));
    InMux I__5773 (
            .O(N__33622),
            .I(N__33616));
    Odrv4 I__5772 (
            .O(N__33619),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_13));
    LocalMux I__5771 (
            .O(N__33616),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_13));
    InMux I__5770 (
            .O(N__33611),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ));
    InMux I__5769 (
            .O(N__33608),
            .I(N__33605));
    LocalMux I__5768 (
            .O(N__33605),
            .I(N__33601));
    InMux I__5767 (
            .O(N__33604),
            .I(N__33598));
    Odrv4 I__5766 (
            .O(N__33601),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_14));
    LocalMux I__5765 (
            .O(N__33598),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_14));
    InMux I__5764 (
            .O(N__33593),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ));
    InMux I__5763 (
            .O(N__33590),
            .I(N__33587));
    LocalMux I__5762 (
            .O(N__33587),
            .I(N__33583));
    InMux I__5761 (
            .O(N__33586),
            .I(N__33580));
    Odrv4 I__5760 (
            .O(N__33583),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_15));
    LocalMux I__5759 (
            .O(N__33580),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_15));
    InMux I__5758 (
            .O(N__33575),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ));
    InMux I__5757 (
            .O(N__33572),
            .I(bfn_12_9_0_));
    InMux I__5756 (
            .O(N__33569),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ));
    InMux I__5755 (
            .O(N__33566),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ));
    InMux I__5754 (
            .O(N__33563),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ));
    InMux I__5753 (
            .O(N__33560),
            .I(N__33556));
    InMux I__5752 (
            .O(N__33559),
            .I(N__33553));
    LocalMux I__5751 (
            .O(N__33556),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_20));
    LocalMux I__5750 (
            .O(N__33553),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_20));
    InMux I__5749 (
            .O(N__33548),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ));
    InMux I__5748 (
            .O(N__33545),
            .I(N__33542));
    LocalMux I__5747 (
            .O(N__33542),
            .I(N__33538));
    InMux I__5746 (
            .O(N__33541),
            .I(N__33535));
    Odrv4 I__5745 (
            .O(N__33538),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_21));
    LocalMux I__5744 (
            .O(N__33535),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_21));
    InMux I__5743 (
            .O(N__33530),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ));
    InMux I__5742 (
            .O(N__33527),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ));
    InMux I__5741 (
            .O(N__33524),
            .I(N__33521));
    LocalMux I__5740 (
            .O(N__33521),
            .I(N__33517));
    InMux I__5739 (
            .O(N__33520),
            .I(N__33514));
    Odrv4 I__5738 (
            .O(N__33517),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_5));
    LocalMux I__5737 (
            .O(N__33514),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_5));
    InMux I__5736 (
            .O(N__33509),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ));
    InMux I__5735 (
            .O(N__33506),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ));
    InMux I__5734 (
            .O(N__33503),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ));
    InMux I__5733 (
            .O(N__33500),
            .I(N__33497));
    LocalMux I__5732 (
            .O(N__33497),
            .I(N__33493));
    InMux I__5731 (
            .O(N__33496),
            .I(N__33490));
    Odrv4 I__5730 (
            .O(N__33493),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_8));
    LocalMux I__5729 (
            .O(N__33490),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_8));
    InMux I__5728 (
            .O(N__33485),
            .I(bfn_12_8_0_));
    InMux I__5727 (
            .O(N__33482),
            .I(N__33479));
    LocalMux I__5726 (
            .O(N__33479),
            .I(N__33475));
    InMux I__5725 (
            .O(N__33478),
            .I(N__33472));
    Odrv4 I__5724 (
            .O(N__33475),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_9));
    LocalMux I__5723 (
            .O(N__33472),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_9));
    InMux I__5722 (
            .O(N__33467),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ));
    InMux I__5721 (
            .O(N__33464),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ));
    InMux I__5720 (
            .O(N__33461),
            .I(N__33457));
    InMux I__5719 (
            .O(N__33460),
            .I(N__33454));
    LocalMux I__5718 (
            .O(N__33457),
            .I(N__33451));
    LocalMux I__5717 (
            .O(N__33454),
            .I(N__33448));
    Odrv4 I__5716 (
            .O(N__33451),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_11));
    Odrv4 I__5715 (
            .O(N__33448),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_11));
    InMux I__5714 (
            .O(N__33443),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ));
    InMux I__5713 (
            .O(N__33440),
            .I(N__33437));
    LocalMux I__5712 (
            .O(N__33437),
            .I(N__33433));
    InMux I__5711 (
            .O(N__33436),
            .I(N__33430));
    Odrv4 I__5710 (
            .O(N__33433),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_12));
    LocalMux I__5709 (
            .O(N__33430),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_12));
    InMux I__5708 (
            .O(N__33425),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ));
    InMux I__5707 (
            .O(N__33422),
            .I(N__33419));
    LocalMux I__5706 (
            .O(N__33419),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ));
    InMux I__5705 (
            .O(N__33416),
            .I(N__33413));
    LocalMux I__5704 (
            .O(N__33413),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ));
    InMux I__5703 (
            .O(N__33410),
            .I(N__33407));
    LocalMux I__5702 (
            .O(N__33407),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ));
    CascadeMux I__5701 (
            .O(N__33404),
            .I(N__33401));
    InMux I__5700 (
            .O(N__33401),
            .I(N__33398));
    LocalMux I__5699 (
            .O(N__33398),
            .I(N__33395));
    Span4Mux_h I__5698 (
            .O(N__33395),
            .I(N__33392));
    Odrv4 I__5697 (
            .O(N__33392),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ));
    CascadeMux I__5696 (
            .O(N__33389),
            .I(N__33386));
    InMux I__5695 (
            .O(N__33386),
            .I(N__33383));
    LocalMux I__5694 (
            .O(N__33383),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ));
    CEMux I__5693 (
            .O(N__33380),
            .I(N__33377));
    LocalMux I__5692 (
            .O(N__33377),
            .I(N__33371));
    CEMux I__5691 (
            .O(N__33376),
            .I(N__33368));
    CEMux I__5690 (
            .O(N__33375),
            .I(N__33364));
    CEMux I__5689 (
            .O(N__33374),
            .I(N__33361));
    Span4Mux_h I__5688 (
            .O(N__33371),
            .I(N__33356));
    LocalMux I__5687 (
            .O(N__33368),
            .I(N__33356));
    CEMux I__5686 (
            .O(N__33367),
            .I(N__33353));
    LocalMux I__5685 (
            .O(N__33364),
            .I(N__33349));
    LocalMux I__5684 (
            .O(N__33361),
            .I(N__33346));
    Span4Mux_v I__5683 (
            .O(N__33356),
            .I(N__33341));
    LocalMux I__5682 (
            .O(N__33353),
            .I(N__33341));
    CEMux I__5681 (
            .O(N__33352),
            .I(N__33338));
    Span4Mux_v I__5680 (
            .O(N__33349),
            .I(N__33335));
    Span4Mux_v I__5679 (
            .O(N__33346),
            .I(N__33332));
    Span4Mux_v I__5678 (
            .O(N__33341),
            .I(N__33329));
    LocalMux I__5677 (
            .O(N__33338),
            .I(N__33326));
    Odrv4 I__5676 (
            .O(N__33335),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__5675 (
            .O(N__33332),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__5674 (
            .O(N__33329),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv12 I__5673 (
            .O(N__33326),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    InMux I__5672 (
            .O(N__33317),
            .I(N__33314));
    LocalMux I__5671 (
            .O(N__33314),
            .I(\phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ));
    InMux I__5670 (
            .O(N__33311),
            .I(N__33308));
    LocalMux I__5669 (
            .O(N__33308),
            .I(N__33304));
    InMux I__5668 (
            .O(N__33307),
            .I(N__33301));
    Span4Mux_h I__5667 (
            .O(N__33304),
            .I(N__33298));
    LocalMux I__5666 (
            .O(N__33301),
            .I(N__33295));
    Odrv4 I__5665 (
            .O(N__33298),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_1));
    Odrv4 I__5664 (
            .O(N__33295),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_1));
    InMux I__5663 (
            .O(N__33290),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ));
    InMux I__5662 (
            .O(N__33287),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ));
    InMux I__5661 (
            .O(N__33284),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ));
    InMux I__5660 (
            .O(N__33281),
            .I(N__33278));
    LocalMux I__5659 (
            .O(N__33278),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ));
    CascadeMux I__5658 (
            .O(N__33275),
            .I(N__33272));
    InMux I__5657 (
            .O(N__33272),
            .I(N__33269));
    LocalMux I__5656 (
            .O(N__33269),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ));
    InMux I__5655 (
            .O(N__33266),
            .I(N__33263));
    LocalMux I__5654 (
            .O(N__33263),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ));
    CascadeMux I__5653 (
            .O(N__33260),
            .I(N__33257));
    InMux I__5652 (
            .O(N__33257),
            .I(N__33254));
    LocalMux I__5651 (
            .O(N__33254),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ));
    CascadeMux I__5650 (
            .O(N__33251),
            .I(N__33248));
    InMux I__5649 (
            .O(N__33248),
            .I(N__33245));
    LocalMux I__5648 (
            .O(N__33245),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ));
    CascadeMux I__5647 (
            .O(N__33242),
            .I(N__33239));
    InMux I__5646 (
            .O(N__33239),
            .I(N__33236));
    LocalMux I__5645 (
            .O(N__33236),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ));
    InMux I__5644 (
            .O(N__33233),
            .I(N__33230));
    LocalMux I__5643 (
            .O(N__33230),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ));
    InMux I__5642 (
            .O(N__33227),
            .I(N__33221));
    InMux I__5641 (
            .O(N__33226),
            .I(N__33221));
    LocalMux I__5640 (
            .O(N__33221),
            .I(N__33218));
    Odrv4 I__5639 (
            .O(N__33218),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ));
    InMux I__5638 (
            .O(N__33215),
            .I(N__33212));
    LocalMux I__5637 (
            .O(N__33212),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ));
    InMux I__5636 (
            .O(N__33209),
            .I(N__33206));
    LocalMux I__5635 (
            .O(N__33206),
            .I(N__33203));
    Span4Mux_v I__5634 (
            .O(N__33203),
            .I(N__33199));
    InMux I__5633 (
            .O(N__33202),
            .I(N__33196));
    Odrv4 I__5632 (
            .O(N__33199),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    LocalMux I__5631 (
            .O(N__33196),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__5630 (
            .O(N__33191),
            .I(bfn_11_23_0_));
    InMux I__5629 (
            .O(N__33188),
            .I(N__33185));
    LocalMux I__5628 (
            .O(N__33185),
            .I(N__33181));
    CascadeMux I__5627 (
            .O(N__33184),
            .I(N__33178));
    Span4Mux_v I__5626 (
            .O(N__33181),
            .I(N__33175));
    InMux I__5625 (
            .O(N__33178),
            .I(N__33172));
    Odrv4 I__5624 (
            .O(N__33175),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    LocalMux I__5623 (
            .O(N__33172),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__5622 (
            .O(N__33167),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__5621 (
            .O(N__33164),
            .I(N__33161));
    LocalMux I__5620 (
            .O(N__33161),
            .I(N__33158));
    Span4Mux_v I__5619 (
            .O(N__33158),
            .I(N__33154));
    InMux I__5618 (
            .O(N__33157),
            .I(N__33151));
    Odrv4 I__5617 (
            .O(N__33154),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    LocalMux I__5616 (
            .O(N__33151),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__5615 (
            .O(N__33146),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__5614 (
            .O(N__33143),
            .I(N__33140));
    LocalMux I__5613 (
            .O(N__33140),
            .I(N__33137));
    Span4Mux_v I__5612 (
            .O(N__33137),
            .I(N__33134));
    Span4Mux_v I__5611 (
            .O(N__33134),
            .I(N__33130));
    InMux I__5610 (
            .O(N__33133),
            .I(N__33127));
    Odrv4 I__5609 (
            .O(N__33130),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    LocalMux I__5608 (
            .O(N__33127),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__5607 (
            .O(N__33122),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__5606 (
            .O(N__33119),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__5605 (
            .O(N__33116),
            .I(N__33113));
    LocalMux I__5604 (
            .O(N__33113),
            .I(N__33109));
    InMux I__5603 (
            .O(N__33112),
            .I(N__33106));
    Span4Mux_v I__5602 (
            .O(N__33109),
            .I(N__33103));
    LocalMux I__5601 (
            .O(N__33106),
            .I(N__33100));
    Span4Mux_h I__5600 (
            .O(N__33103),
            .I(N__33095));
    Span4Mux_v I__5599 (
            .O(N__33100),
            .I(N__33095));
    Span4Mux_v I__5598 (
            .O(N__33095),
            .I(N__33092));
    Odrv4 I__5597 (
            .O(N__33092),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__5596 (
            .O(N__33089),
            .I(N__33086));
    LocalMux I__5595 (
            .O(N__33086),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ));
    InMux I__5594 (
            .O(N__33083),
            .I(N__33080));
    LocalMux I__5593 (
            .O(N__33080),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ));
    CascadeMux I__5592 (
            .O(N__33077),
            .I(N__33074));
    InMux I__5591 (
            .O(N__33074),
            .I(N__33071));
    LocalMux I__5590 (
            .O(N__33071),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ));
    InMux I__5589 (
            .O(N__33068),
            .I(N__33065));
    LocalMux I__5588 (
            .O(N__33065),
            .I(N__33062));
    Span4Mux_v I__5587 (
            .O(N__33062),
            .I(N__33058));
    InMux I__5586 (
            .O(N__33061),
            .I(N__33055));
    Odrv4 I__5585 (
            .O(N__33058),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__5584 (
            .O(N__33055),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__5583 (
            .O(N__33050),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__5582 (
            .O(N__33047),
            .I(N__33041));
    InMux I__5581 (
            .O(N__33046),
            .I(N__33041));
    LocalMux I__5580 (
            .O(N__33041),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__5579 (
            .O(N__33038),
            .I(bfn_11_22_0_));
    InMux I__5578 (
            .O(N__33035),
            .I(N__33032));
    LocalMux I__5577 (
            .O(N__33032),
            .I(N__33029));
    Span4Mux_h I__5576 (
            .O(N__33029),
            .I(N__33026));
    Span4Mux_v I__5575 (
            .O(N__33026),
            .I(N__33022));
    InMux I__5574 (
            .O(N__33025),
            .I(N__33019));
    Odrv4 I__5573 (
            .O(N__33022),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__5572 (
            .O(N__33019),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__5571 (
            .O(N__33014),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__5570 (
            .O(N__33011),
            .I(N__33008));
    LocalMux I__5569 (
            .O(N__33008),
            .I(N__33005));
    Span4Mux_v I__5568 (
            .O(N__33005),
            .I(N__33002));
    Span4Mux_v I__5567 (
            .O(N__33002),
            .I(N__32998));
    InMux I__5566 (
            .O(N__33001),
            .I(N__32995));
    Odrv4 I__5565 (
            .O(N__32998),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__5564 (
            .O(N__32995),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__5563 (
            .O(N__32990),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__5562 (
            .O(N__32987),
            .I(N__32984));
    LocalMux I__5561 (
            .O(N__32984),
            .I(N__32980));
    CascadeMux I__5560 (
            .O(N__32983),
            .I(N__32977));
    Span4Mux_v I__5559 (
            .O(N__32980),
            .I(N__32974));
    InMux I__5558 (
            .O(N__32977),
            .I(N__32971));
    Odrv4 I__5557 (
            .O(N__32974),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    LocalMux I__5556 (
            .O(N__32971),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__5555 (
            .O(N__32966),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__5554 (
            .O(N__32963),
            .I(N__32960));
    LocalMux I__5553 (
            .O(N__32960),
            .I(N__32957));
    Span4Mux_h I__5552 (
            .O(N__32957),
            .I(N__32954));
    Span4Mux_v I__5551 (
            .O(N__32954),
            .I(N__32951));
    Span4Mux_v I__5550 (
            .O(N__32951),
            .I(N__32947));
    InMux I__5549 (
            .O(N__32950),
            .I(N__32944));
    Odrv4 I__5548 (
            .O(N__32947),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__5547 (
            .O(N__32944),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__5546 (
            .O(N__32939),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__5545 (
            .O(N__32936),
            .I(N__32933));
    LocalMux I__5544 (
            .O(N__32933),
            .I(N__32929));
    CascadeMux I__5543 (
            .O(N__32932),
            .I(N__32926));
    Span12Mux_v I__5542 (
            .O(N__32929),
            .I(N__32923));
    InMux I__5541 (
            .O(N__32926),
            .I(N__32920));
    Odrv12 I__5540 (
            .O(N__32923),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__5539 (
            .O(N__32920),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__5538 (
            .O(N__32915),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__5537 (
            .O(N__32912),
            .I(N__32909));
    LocalMux I__5536 (
            .O(N__32909),
            .I(N__32906));
    Span4Mux_v I__5535 (
            .O(N__32906),
            .I(N__32902));
    InMux I__5534 (
            .O(N__32905),
            .I(N__32899));
    Odrv4 I__5533 (
            .O(N__32902),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__5532 (
            .O(N__32899),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__5531 (
            .O(N__32894),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__5530 (
            .O(N__32891),
            .I(N__32888));
    LocalMux I__5529 (
            .O(N__32888),
            .I(N__32885));
    Span4Mux_v I__5528 (
            .O(N__32885),
            .I(N__32881));
    InMux I__5527 (
            .O(N__32884),
            .I(N__32878));
    Odrv4 I__5526 (
            .O(N__32881),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    LocalMux I__5525 (
            .O(N__32878),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__5524 (
            .O(N__32873),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__5523 (
            .O(N__32870),
            .I(N__32867));
    LocalMux I__5522 (
            .O(N__32867),
            .I(N__32864));
    Span4Mux_v I__5521 (
            .O(N__32864),
            .I(N__32860));
    InMux I__5520 (
            .O(N__32863),
            .I(N__32857));
    Odrv4 I__5519 (
            .O(N__32860),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__5518 (
            .O(N__32857),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__5517 (
            .O(N__32852),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__5516 (
            .O(N__32849),
            .I(N__32846));
    LocalMux I__5515 (
            .O(N__32846),
            .I(N__32843));
    Span4Mux_h I__5514 (
            .O(N__32843),
            .I(N__32840));
    Span4Mux_v I__5513 (
            .O(N__32840),
            .I(N__32836));
    InMux I__5512 (
            .O(N__32839),
            .I(N__32833));
    Odrv4 I__5511 (
            .O(N__32836),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__5510 (
            .O(N__32833),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__5509 (
            .O(N__32828),
            .I(bfn_11_21_0_));
    InMux I__5508 (
            .O(N__32825),
            .I(N__32822));
    LocalMux I__5507 (
            .O(N__32822),
            .I(N__32819));
    Span4Mux_v I__5506 (
            .O(N__32819),
            .I(N__32815));
    InMux I__5505 (
            .O(N__32818),
            .I(N__32812));
    Odrv4 I__5504 (
            .O(N__32815),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    LocalMux I__5503 (
            .O(N__32812),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__5502 (
            .O(N__32807),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__5501 (
            .O(N__32804),
            .I(N__32801));
    LocalMux I__5500 (
            .O(N__32801),
            .I(N__32798));
    Span4Mux_h I__5499 (
            .O(N__32798),
            .I(N__32795));
    Span4Mux_v I__5498 (
            .O(N__32795),
            .I(N__32792));
    Span4Mux_v I__5497 (
            .O(N__32792),
            .I(N__32788));
    InMux I__5496 (
            .O(N__32791),
            .I(N__32785));
    Odrv4 I__5495 (
            .O(N__32788),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__5494 (
            .O(N__32785),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__5493 (
            .O(N__32780),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__5492 (
            .O(N__32777),
            .I(N__32774));
    LocalMux I__5491 (
            .O(N__32774),
            .I(N__32771));
    Span4Mux_h I__5490 (
            .O(N__32771),
            .I(N__32768));
    Span4Mux_v I__5489 (
            .O(N__32768),
            .I(N__32764));
    InMux I__5488 (
            .O(N__32767),
            .I(N__32761));
    Odrv4 I__5487 (
            .O(N__32764),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    LocalMux I__5486 (
            .O(N__32761),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__5485 (
            .O(N__32756),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__5484 (
            .O(N__32753),
            .I(N__32750));
    LocalMux I__5483 (
            .O(N__32750),
            .I(N__32747));
    Span4Mux_h I__5482 (
            .O(N__32747),
            .I(N__32744));
    Span4Mux_v I__5481 (
            .O(N__32744),
            .I(N__32740));
    InMux I__5480 (
            .O(N__32743),
            .I(N__32737));
    Odrv4 I__5479 (
            .O(N__32740),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    LocalMux I__5478 (
            .O(N__32737),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__5477 (
            .O(N__32732),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__5476 (
            .O(N__32729),
            .I(N__32726));
    LocalMux I__5475 (
            .O(N__32726),
            .I(N__32722));
    CascadeMux I__5474 (
            .O(N__32725),
            .I(N__32719));
    Span4Mux_v I__5473 (
            .O(N__32722),
            .I(N__32716));
    InMux I__5472 (
            .O(N__32719),
            .I(N__32713));
    Odrv4 I__5471 (
            .O(N__32716),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__5470 (
            .O(N__32713),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__5469 (
            .O(N__32708),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__5468 (
            .O(N__32705),
            .I(N__32702));
    LocalMux I__5467 (
            .O(N__32702),
            .I(N__32699));
    Span4Mux_v I__5466 (
            .O(N__32699),
            .I(N__32695));
    InMux I__5465 (
            .O(N__32698),
            .I(N__32692));
    Odrv4 I__5464 (
            .O(N__32695),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__5463 (
            .O(N__32692),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__5462 (
            .O(N__32687),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__5461 (
            .O(N__32684),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_29 ));
    InMux I__5460 (
            .O(N__32681),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_30 ));
    CEMux I__5459 (
            .O(N__32678),
            .I(N__32672));
    CEMux I__5458 (
            .O(N__32677),
            .I(N__32669));
    CEMux I__5457 (
            .O(N__32676),
            .I(N__32666));
    CEMux I__5456 (
            .O(N__32675),
            .I(N__32663));
    LocalMux I__5455 (
            .O(N__32672),
            .I(N__32660));
    LocalMux I__5454 (
            .O(N__32669),
            .I(N__32655));
    LocalMux I__5453 (
            .O(N__32666),
            .I(N__32655));
    LocalMux I__5452 (
            .O(N__32663),
            .I(N__32652));
    Span4Mux_v I__5451 (
            .O(N__32660),
            .I(N__32647));
    Span4Mux_v I__5450 (
            .O(N__32655),
            .I(N__32647));
    Span12Mux_h I__5449 (
            .O(N__32652),
            .I(N__32644));
    Odrv4 I__5448 (
            .O(N__32647),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv12 I__5447 (
            .O(N__32644),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    InMux I__5446 (
            .O(N__32639),
            .I(N__32633));
    InMux I__5445 (
            .O(N__32638),
            .I(N__32633));
    LocalMux I__5444 (
            .O(N__32633),
            .I(N__32630));
    Span4Mux_h I__5443 (
            .O(N__32630),
            .I(N__32627));
    Span4Mux_v I__5442 (
            .O(N__32627),
            .I(N__32624));
    Odrv4 I__5441 (
            .O(N__32624),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    CascadeMux I__5440 (
            .O(N__32621),
            .I(N__32618));
    InMux I__5439 (
            .O(N__32618),
            .I(N__32614));
    InMux I__5438 (
            .O(N__32617),
            .I(N__32611));
    LocalMux I__5437 (
            .O(N__32614),
            .I(N__32608));
    LocalMux I__5436 (
            .O(N__32611),
            .I(N__32603));
    Span4Mux_h I__5435 (
            .O(N__32608),
            .I(N__32603));
    Span4Mux_v I__5434 (
            .O(N__32603),
            .I(N__32600));
    Odrv4 I__5433 (
            .O(N__32600),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__5432 (
            .O(N__32597),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__5431 (
            .O(N__32594),
            .I(N__32591));
    LocalMux I__5430 (
            .O(N__32591),
            .I(N__32588));
    Span4Mux_v I__5429 (
            .O(N__32588),
            .I(N__32584));
    InMux I__5428 (
            .O(N__32587),
            .I(N__32581));
    Odrv4 I__5427 (
            .O(N__32584),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__5426 (
            .O(N__32581),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__5425 (
            .O(N__32576),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__5424 (
            .O(N__32573),
            .I(N__32570));
    LocalMux I__5423 (
            .O(N__32570),
            .I(N__32567));
    Span4Mux_v I__5422 (
            .O(N__32567),
            .I(N__32563));
    InMux I__5421 (
            .O(N__32566),
            .I(N__32560));
    Odrv4 I__5420 (
            .O(N__32563),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    LocalMux I__5419 (
            .O(N__32560),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__5418 (
            .O(N__32555),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__5417 (
            .O(N__32552),
            .I(N__32549));
    LocalMux I__5416 (
            .O(N__32549),
            .I(N__32545));
    InMux I__5415 (
            .O(N__32548),
            .I(N__32542));
    Span4Mux_h I__5414 (
            .O(N__32545),
            .I(N__32537));
    LocalMux I__5413 (
            .O(N__32542),
            .I(N__32537));
    Span4Mux_v I__5412 (
            .O(N__32537),
            .I(N__32534));
    Odrv4 I__5411 (
            .O(N__32534),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__5410 (
            .O(N__32531),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__5409 (
            .O(N__32528),
            .I(N__32524));
    InMux I__5408 (
            .O(N__32527),
            .I(N__32519));
    InMux I__5407 (
            .O(N__32524),
            .I(N__32519));
    LocalMux I__5406 (
            .O(N__32519),
            .I(N__32516));
    Span12Mux_v I__5405 (
            .O(N__32516),
            .I(N__32513));
    Odrv12 I__5404 (
            .O(N__32513),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__5403 (
            .O(N__32510),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__5402 (
            .O(N__32507),
            .I(N__32504));
    LocalMux I__5401 (
            .O(N__32504),
            .I(N__32500));
    CascadeMux I__5400 (
            .O(N__32503),
            .I(N__32497));
    Span4Mux_v I__5399 (
            .O(N__32500),
            .I(N__32494));
    InMux I__5398 (
            .O(N__32497),
            .I(N__32491));
    Odrv4 I__5397 (
            .O(N__32494),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    LocalMux I__5396 (
            .O(N__32491),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__5395 (
            .O(N__32486),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__5394 (
            .O(N__32483),
            .I(N__32479));
    CascadeMux I__5393 (
            .O(N__32482),
            .I(N__32476));
    InMux I__5392 (
            .O(N__32479),
            .I(N__32471));
    InMux I__5391 (
            .O(N__32476),
            .I(N__32471));
    LocalMux I__5390 (
            .O(N__32471),
            .I(N__32467));
    InMux I__5389 (
            .O(N__32470),
            .I(N__32464));
    Span12Mux_s11_v I__5388 (
            .O(N__32467),
            .I(N__32461));
    LocalMux I__5387 (
            .O(N__32464),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ));
    Odrv12 I__5386 (
            .O(N__32461),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ));
    InMux I__5385 (
            .O(N__32456),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_21 ));
    InMux I__5384 (
            .O(N__32453),
            .I(N__32447));
    InMux I__5383 (
            .O(N__32452),
            .I(N__32447));
    LocalMux I__5382 (
            .O(N__32447),
            .I(N__32443));
    InMux I__5381 (
            .O(N__32446),
            .I(N__32440));
    Span12Mux_v I__5380 (
            .O(N__32443),
            .I(N__32437));
    LocalMux I__5379 (
            .O(N__32440),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ));
    Odrv12 I__5378 (
            .O(N__32437),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ));
    InMux I__5377 (
            .O(N__32432),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_22 ));
    CascadeMux I__5376 (
            .O(N__32429),
            .I(N__32425));
    CascadeMux I__5375 (
            .O(N__32428),
            .I(N__32422));
    InMux I__5374 (
            .O(N__32425),
            .I(N__32417));
    InMux I__5373 (
            .O(N__32422),
            .I(N__32417));
    LocalMux I__5372 (
            .O(N__32417),
            .I(N__32413));
    InMux I__5371 (
            .O(N__32416),
            .I(N__32410));
    Span12Mux_v I__5370 (
            .O(N__32413),
            .I(N__32407));
    LocalMux I__5369 (
            .O(N__32410),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ));
    Odrv12 I__5368 (
            .O(N__32407),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ));
    InMux I__5367 (
            .O(N__32402),
            .I(bfn_11_19_0_));
    InMux I__5366 (
            .O(N__32399),
            .I(N__32393));
    InMux I__5365 (
            .O(N__32398),
            .I(N__32393));
    LocalMux I__5364 (
            .O(N__32393),
            .I(N__32389));
    InMux I__5363 (
            .O(N__32392),
            .I(N__32386));
    Span12Mux_v I__5362 (
            .O(N__32389),
            .I(N__32383));
    LocalMux I__5361 (
            .O(N__32386),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ));
    Odrv12 I__5360 (
            .O(N__32383),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ));
    InMux I__5359 (
            .O(N__32378),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_24 ));
    CascadeMux I__5358 (
            .O(N__32375),
            .I(N__32371));
    CascadeMux I__5357 (
            .O(N__32374),
            .I(N__32368));
    InMux I__5356 (
            .O(N__32371),
            .I(N__32362));
    InMux I__5355 (
            .O(N__32368),
            .I(N__32362));
    InMux I__5354 (
            .O(N__32367),
            .I(N__32359));
    LocalMux I__5353 (
            .O(N__32362),
            .I(N__32356));
    LocalMux I__5352 (
            .O(N__32359),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ));
    Odrv12 I__5351 (
            .O(N__32356),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ));
    InMux I__5350 (
            .O(N__32351),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_25 ));
    InMux I__5349 (
            .O(N__32348),
            .I(N__32341));
    InMux I__5348 (
            .O(N__32347),
            .I(N__32341));
    InMux I__5347 (
            .O(N__32346),
            .I(N__32338));
    LocalMux I__5346 (
            .O(N__32341),
            .I(N__32335));
    LocalMux I__5345 (
            .O(N__32338),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ));
    Odrv12 I__5344 (
            .O(N__32335),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ));
    InMux I__5343 (
            .O(N__32330),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_26 ));
    InMux I__5342 (
            .O(N__32327),
            .I(N__32321));
    InMux I__5341 (
            .O(N__32326),
            .I(N__32321));
    LocalMux I__5340 (
            .O(N__32321),
            .I(N__32317));
    InMux I__5339 (
            .O(N__32320),
            .I(N__32314));
    Span4Mux_h I__5338 (
            .O(N__32317),
            .I(N__32311));
    LocalMux I__5337 (
            .O(N__32314),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ));
    Odrv4 I__5336 (
            .O(N__32311),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ));
    InMux I__5335 (
            .O(N__32306),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_27 ));
    InMux I__5334 (
            .O(N__32303),
            .I(N__32297));
    InMux I__5333 (
            .O(N__32302),
            .I(N__32297));
    LocalMux I__5332 (
            .O(N__32297),
            .I(N__32293));
    InMux I__5331 (
            .O(N__32296),
            .I(N__32290));
    Span4Mux_v I__5330 (
            .O(N__32293),
            .I(N__32287));
    LocalMux I__5329 (
            .O(N__32290),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ));
    Odrv4 I__5328 (
            .O(N__32287),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ));
    InMux I__5327 (
            .O(N__32282),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_28 ));
    InMux I__5326 (
            .O(N__32279),
            .I(N__32276));
    LocalMux I__5325 (
            .O(N__32276),
            .I(N__32272));
    InMux I__5324 (
            .O(N__32275),
            .I(N__32269));
    Span4Mux_v I__5323 (
            .O(N__32272),
            .I(N__32266));
    LocalMux I__5322 (
            .O(N__32269),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ));
    Odrv4 I__5321 (
            .O(N__32266),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ));
    InMux I__5320 (
            .O(N__32261),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_12 ));
    InMux I__5319 (
            .O(N__32258),
            .I(N__32254));
    InMux I__5318 (
            .O(N__32257),
            .I(N__32251));
    LocalMux I__5317 (
            .O(N__32254),
            .I(N__32248));
    LocalMux I__5316 (
            .O(N__32251),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ));
    Odrv12 I__5315 (
            .O(N__32248),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ));
    InMux I__5314 (
            .O(N__32243),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_13 ));
    InMux I__5313 (
            .O(N__32240),
            .I(N__32236));
    InMux I__5312 (
            .O(N__32239),
            .I(N__32233));
    LocalMux I__5311 (
            .O(N__32236),
            .I(N__32230));
    LocalMux I__5310 (
            .O(N__32233),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ));
    Odrv12 I__5309 (
            .O(N__32230),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ));
    InMux I__5308 (
            .O(N__32225),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_14 ));
    InMux I__5307 (
            .O(N__32222),
            .I(bfn_11_18_0_));
    InMux I__5306 (
            .O(N__32219),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_16 ));
    InMux I__5305 (
            .O(N__32216),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_17 ));
    InMux I__5304 (
            .O(N__32213),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_18 ));
    CascadeMux I__5303 (
            .O(N__32210),
            .I(N__32206));
    CascadeMux I__5302 (
            .O(N__32209),
            .I(N__32203));
    InMux I__5301 (
            .O(N__32206),
            .I(N__32198));
    InMux I__5300 (
            .O(N__32203),
            .I(N__32198));
    LocalMux I__5299 (
            .O(N__32198),
            .I(N__32194));
    InMux I__5298 (
            .O(N__32197),
            .I(N__32191));
    Sp12to4 I__5297 (
            .O(N__32194),
            .I(N__32188));
    LocalMux I__5296 (
            .O(N__32191),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ));
    Odrv12 I__5295 (
            .O(N__32188),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ));
    InMux I__5294 (
            .O(N__32183),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_19 ));
    InMux I__5293 (
            .O(N__32180),
            .I(N__32174));
    InMux I__5292 (
            .O(N__32179),
            .I(N__32174));
    LocalMux I__5291 (
            .O(N__32174),
            .I(N__32171));
    Span4Mux_h I__5290 (
            .O(N__32171),
            .I(N__32167));
    InMux I__5289 (
            .O(N__32170),
            .I(N__32164));
    Span4Mux_v I__5288 (
            .O(N__32167),
            .I(N__32161));
    LocalMux I__5287 (
            .O(N__32164),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ));
    Odrv4 I__5286 (
            .O(N__32161),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ));
    InMux I__5285 (
            .O(N__32156),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_20 ));
    InMux I__5284 (
            .O(N__32153),
            .I(N__32149));
    InMux I__5283 (
            .O(N__32152),
            .I(N__32146));
    LocalMux I__5282 (
            .O(N__32149),
            .I(N__32143));
    LocalMux I__5281 (
            .O(N__32146),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ));
    Odrv12 I__5280 (
            .O(N__32143),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ));
    InMux I__5279 (
            .O(N__32138),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_4 ));
    InMux I__5278 (
            .O(N__32135),
            .I(N__32132));
    LocalMux I__5277 (
            .O(N__32132),
            .I(N__32128));
    InMux I__5276 (
            .O(N__32131),
            .I(N__32125));
    Span4Mux_v I__5275 (
            .O(N__32128),
            .I(N__32122));
    LocalMux I__5274 (
            .O(N__32125),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ));
    Odrv4 I__5273 (
            .O(N__32122),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ));
    InMux I__5272 (
            .O(N__32117),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_5 ));
    InMux I__5271 (
            .O(N__32114),
            .I(N__32110));
    InMux I__5270 (
            .O(N__32113),
            .I(N__32107));
    LocalMux I__5269 (
            .O(N__32110),
            .I(N__32104));
    LocalMux I__5268 (
            .O(N__32107),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ));
    Odrv12 I__5267 (
            .O(N__32104),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ));
    InMux I__5266 (
            .O(N__32099),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_6 ));
    InMux I__5265 (
            .O(N__32096),
            .I(N__32092));
    InMux I__5264 (
            .O(N__32095),
            .I(N__32089));
    LocalMux I__5263 (
            .O(N__32092),
            .I(N__32086));
    LocalMux I__5262 (
            .O(N__32089),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ));
    Odrv12 I__5261 (
            .O(N__32086),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ));
    InMux I__5260 (
            .O(N__32081),
            .I(bfn_11_17_0_));
    InMux I__5259 (
            .O(N__32078),
            .I(N__32074));
    InMux I__5258 (
            .O(N__32077),
            .I(N__32071));
    LocalMux I__5257 (
            .O(N__32074),
            .I(N__32068));
    LocalMux I__5256 (
            .O(N__32071),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ));
    Odrv12 I__5255 (
            .O(N__32068),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ));
    InMux I__5254 (
            .O(N__32063),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_8 ));
    InMux I__5253 (
            .O(N__32060),
            .I(N__32057));
    LocalMux I__5252 (
            .O(N__32057),
            .I(N__32053));
    InMux I__5251 (
            .O(N__32056),
            .I(N__32050));
    Span4Mux_h I__5250 (
            .O(N__32053),
            .I(N__32047));
    LocalMux I__5249 (
            .O(N__32050),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ));
    Odrv4 I__5248 (
            .O(N__32047),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ));
    InMux I__5247 (
            .O(N__32042),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_9 ));
    InMux I__5246 (
            .O(N__32039),
            .I(N__32035));
    InMux I__5245 (
            .O(N__32038),
            .I(N__32032));
    LocalMux I__5244 (
            .O(N__32035),
            .I(N__32029));
    LocalMux I__5243 (
            .O(N__32032),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ));
    Odrv12 I__5242 (
            .O(N__32029),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ));
    InMux I__5241 (
            .O(N__32024),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_10 ));
    InMux I__5240 (
            .O(N__32021),
            .I(N__32018));
    LocalMux I__5239 (
            .O(N__32018),
            .I(N__32014));
    InMux I__5238 (
            .O(N__32017),
            .I(N__32011));
    Span4Mux_h I__5237 (
            .O(N__32014),
            .I(N__32008));
    LocalMux I__5236 (
            .O(N__32011),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ));
    Odrv4 I__5235 (
            .O(N__32008),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ));
    InMux I__5234 (
            .O(N__32003),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_11 ));
    CascadeMux I__5233 (
            .O(N__32000),
            .I(N__31997));
    InMux I__5232 (
            .O(N__31997),
            .I(N__31994));
    LocalMux I__5231 (
            .O(N__31994),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ));
    InMux I__5230 (
            .O(N__31991),
            .I(N__31988));
    LocalMux I__5229 (
            .O(N__31988),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ));
    InMux I__5228 (
            .O(N__31985),
            .I(N__31982));
    LocalMux I__5227 (
            .O(N__31982),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt28 ));
    CascadeMux I__5226 (
            .O(N__31979),
            .I(N__31975));
    InMux I__5225 (
            .O(N__31978),
            .I(N__31972));
    InMux I__5224 (
            .O(N__31975),
            .I(N__31969));
    LocalMux I__5223 (
            .O(N__31972),
            .I(\phase_controller_inst1.stoper_hc.counter ));
    LocalMux I__5222 (
            .O(N__31969),
            .I(\phase_controller_inst1.stoper_hc.counter ));
    InMux I__5221 (
            .O(N__31964),
            .I(N__31961));
    LocalMux I__5220 (
            .O(N__31961),
            .I(N__31957));
    InMux I__5219 (
            .O(N__31960),
            .I(N__31954));
    Span4Mux_v I__5218 (
            .O(N__31957),
            .I(N__31951));
    LocalMux I__5217 (
            .O(N__31954),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ));
    Odrv4 I__5216 (
            .O(N__31951),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ));
    InMux I__5215 (
            .O(N__31946),
            .I(N__31943));
    LocalMux I__5214 (
            .O(N__31943),
            .I(N__31939));
    InMux I__5213 (
            .O(N__31942),
            .I(N__31936));
    Span4Mux_v I__5212 (
            .O(N__31939),
            .I(N__31933));
    LocalMux I__5211 (
            .O(N__31936),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ));
    Odrv4 I__5210 (
            .O(N__31933),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ));
    InMux I__5209 (
            .O(N__31928),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_0 ));
    InMux I__5208 (
            .O(N__31925),
            .I(N__31922));
    LocalMux I__5207 (
            .O(N__31922),
            .I(N__31918));
    InMux I__5206 (
            .O(N__31921),
            .I(N__31915));
    Span4Mux_v I__5205 (
            .O(N__31918),
            .I(N__31912));
    LocalMux I__5204 (
            .O(N__31915),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ));
    Odrv4 I__5203 (
            .O(N__31912),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ));
    InMux I__5202 (
            .O(N__31907),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_1 ));
    InMux I__5201 (
            .O(N__31904),
            .I(N__31900));
    InMux I__5200 (
            .O(N__31903),
            .I(N__31897));
    LocalMux I__5199 (
            .O(N__31900),
            .I(N__31894));
    LocalMux I__5198 (
            .O(N__31897),
            .I(N__31889));
    Span4Mux_v I__5197 (
            .O(N__31894),
            .I(N__31889));
    Odrv4 I__5196 (
            .O(N__31889),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_3 ));
    InMux I__5195 (
            .O(N__31886),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_2 ));
    InMux I__5194 (
            .O(N__31883),
            .I(N__31880));
    LocalMux I__5193 (
            .O(N__31880),
            .I(N__31876));
    InMux I__5192 (
            .O(N__31879),
            .I(N__31873));
    Span4Mux_v I__5191 (
            .O(N__31876),
            .I(N__31870));
    LocalMux I__5190 (
            .O(N__31873),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ));
    Odrv4 I__5189 (
            .O(N__31870),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ));
    InMux I__5188 (
            .O(N__31865),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_3 ));
    InMux I__5187 (
            .O(N__31862),
            .I(N__31859));
    LocalMux I__5186 (
            .O(N__31859),
            .I(N__31856));
    Span4Mux_v I__5185 (
            .O(N__31856),
            .I(N__31853));
    Odrv4 I__5184 (
            .O(N__31853),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt22 ));
    CascadeMux I__5183 (
            .O(N__31850),
            .I(N__31847));
    InMux I__5182 (
            .O(N__31847),
            .I(N__31844));
    LocalMux I__5181 (
            .O(N__31844),
            .I(N__31841));
    Span4Mux_v I__5180 (
            .O(N__31841),
            .I(N__31838));
    Odrv4 I__5179 (
            .O(N__31838),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ));
    InMux I__5178 (
            .O(N__31835),
            .I(N__31832));
    LocalMux I__5177 (
            .O(N__31832),
            .I(N__31829));
    Odrv4 I__5176 (
            .O(N__31829),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ));
    CascadeMux I__5175 (
            .O(N__31826),
            .I(N__31823));
    InMux I__5174 (
            .O(N__31823),
            .I(N__31820));
    LocalMux I__5173 (
            .O(N__31820),
            .I(N__31817));
    Odrv12 I__5172 (
            .O(N__31817),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt24 ));
    InMux I__5171 (
            .O(N__31814),
            .I(N__31811));
    LocalMux I__5170 (
            .O(N__31811),
            .I(N__31808));
    Span4Mux_h I__5169 (
            .O(N__31808),
            .I(N__31805));
    Odrv4 I__5168 (
            .O(N__31805),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt26 ));
    CascadeMux I__5167 (
            .O(N__31802),
            .I(N__31799));
    InMux I__5166 (
            .O(N__31799),
            .I(N__31796));
    LocalMux I__5165 (
            .O(N__31796),
            .I(N__31793));
    Odrv4 I__5164 (
            .O(N__31793),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ));
    InMux I__5163 (
            .O(N__31790),
            .I(bfn_11_15_0_));
    InMux I__5162 (
            .O(N__31787),
            .I(N__31782));
    InMux I__5161 (
            .O(N__31786),
            .I(N__31775));
    InMux I__5160 (
            .O(N__31785),
            .I(N__31763));
    LocalMux I__5159 (
            .O(N__31782),
            .I(N__31760));
    InMux I__5158 (
            .O(N__31781),
            .I(N__31747));
    InMux I__5157 (
            .O(N__31780),
            .I(N__31747));
    InMux I__5156 (
            .O(N__31779),
            .I(N__31747));
    InMux I__5155 (
            .O(N__31778),
            .I(N__31747));
    LocalMux I__5154 (
            .O(N__31775),
            .I(N__31744));
    InMux I__5153 (
            .O(N__31774),
            .I(N__31737));
    InMux I__5152 (
            .O(N__31773),
            .I(N__31737));
    InMux I__5151 (
            .O(N__31772),
            .I(N__31737));
    InMux I__5150 (
            .O(N__31771),
            .I(N__31720));
    InMux I__5149 (
            .O(N__31770),
            .I(N__31720));
    InMux I__5148 (
            .O(N__31769),
            .I(N__31720));
    InMux I__5147 (
            .O(N__31768),
            .I(N__31713));
    InMux I__5146 (
            .O(N__31767),
            .I(N__31713));
    InMux I__5145 (
            .O(N__31766),
            .I(N__31713));
    LocalMux I__5144 (
            .O(N__31763),
            .I(N__31710));
    Span4Mux_h I__5143 (
            .O(N__31760),
            .I(N__31707));
    InMux I__5142 (
            .O(N__31759),
            .I(N__31698));
    InMux I__5141 (
            .O(N__31758),
            .I(N__31698));
    InMux I__5140 (
            .O(N__31757),
            .I(N__31698));
    InMux I__5139 (
            .O(N__31756),
            .I(N__31698));
    LocalMux I__5138 (
            .O(N__31747),
            .I(N__31693));
    Span12Mux_v I__5137 (
            .O(N__31744),
            .I(N__31693));
    LocalMux I__5136 (
            .O(N__31737),
            .I(N__31690));
    InMux I__5135 (
            .O(N__31736),
            .I(N__31685));
    InMux I__5134 (
            .O(N__31735),
            .I(N__31685));
    InMux I__5133 (
            .O(N__31734),
            .I(N__31682));
    InMux I__5132 (
            .O(N__31733),
            .I(N__31677));
    InMux I__5131 (
            .O(N__31732),
            .I(N__31677));
    InMux I__5130 (
            .O(N__31731),
            .I(N__31668));
    InMux I__5129 (
            .O(N__31730),
            .I(N__31668));
    InMux I__5128 (
            .O(N__31729),
            .I(N__31668));
    InMux I__5127 (
            .O(N__31728),
            .I(N__31668));
    InMux I__5126 (
            .O(N__31727),
            .I(N__31665));
    LocalMux I__5125 (
            .O(N__31720),
            .I(N__31660));
    LocalMux I__5124 (
            .O(N__31713),
            .I(N__31660));
    Odrv4 I__5123 (
            .O(N__31710),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5122 (
            .O(N__31707),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5121 (
            .O(N__31698),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__5120 (
            .O(N__31693),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5119 (
            .O(N__31690),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5118 (
            .O(N__31685),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5117 (
            .O(N__31682),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5116 (
            .O(N__31677),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5115 (
            .O(N__31668),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5114 (
            .O(N__31665),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5113 (
            .O(N__31660),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__5112 (
            .O(N__31637),
            .I(N__31634));
    LocalMux I__5111 (
            .O(N__31634),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    CascadeMux I__5110 (
            .O(N__31631),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_));
    InMux I__5109 (
            .O(N__31628),
            .I(N__31625));
    LocalMux I__5108 (
            .O(N__31625),
            .I(N__31622));
    Span4Mux_h I__5107 (
            .O(N__31622),
            .I(N__31619));
    Odrv4 I__5106 (
            .O(N__31619),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ));
    CascadeMux I__5105 (
            .O(N__31616),
            .I(N__31613));
    InMux I__5104 (
            .O(N__31613),
            .I(N__31610));
    LocalMux I__5103 (
            .O(N__31610),
            .I(N__31607));
    Span4Mux_v I__5102 (
            .O(N__31607),
            .I(N__31604));
    Span4Mux_v I__5101 (
            .O(N__31604),
            .I(N__31601));
    Odrv4 I__5100 (
            .O(N__31601),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ));
    InMux I__5099 (
            .O(N__31598),
            .I(N__31595));
    LocalMux I__5098 (
            .O(N__31595),
            .I(\phase_controller_inst1.stoper_hc.counter_i_11 ));
    InMux I__5097 (
            .O(N__31592),
            .I(N__31589));
    LocalMux I__5096 (
            .O(N__31589),
            .I(N__31586));
    Span4Mux_v I__5095 (
            .O(N__31586),
            .I(N__31583));
    Odrv4 I__5094 (
            .O(N__31583),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ));
    CascadeMux I__5093 (
            .O(N__31580),
            .I(N__31577));
    InMux I__5092 (
            .O(N__31577),
            .I(N__31574));
    LocalMux I__5091 (
            .O(N__31574),
            .I(\phase_controller_inst1.stoper_hc.counter_i_12 ));
    InMux I__5090 (
            .O(N__31571),
            .I(N__31568));
    LocalMux I__5089 (
            .O(N__31568),
            .I(N__31565));
    Odrv12 I__5088 (
            .O(N__31565),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ));
    CascadeMux I__5087 (
            .O(N__31562),
            .I(N__31559));
    InMux I__5086 (
            .O(N__31559),
            .I(N__31556));
    LocalMux I__5085 (
            .O(N__31556),
            .I(N__31553));
    Odrv4 I__5084 (
            .O(N__31553),
            .I(\phase_controller_inst1.stoper_hc.counter_i_13 ));
    InMux I__5083 (
            .O(N__31550),
            .I(N__31547));
    LocalMux I__5082 (
            .O(N__31547),
            .I(N__31544));
    Span4Mux_v I__5081 (
            .O(N__31544),
            .I(N__31541));
    Odrv4 I__5080 (
            .O(N__31541),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ));
    CascadeMux I__5079 (
            .O(N__31538),
            .I(N__31535));
    InMux I__5078 (
            .O(N__31535),
            .I(N__31532));
    LocalMux I__5077 (
            .O(N__31532),
            .I(N__31529));
    Odrv4 I__5076 (
            .O(N__31529),
            .I(\phase_controller_inst1.stoper_hc.counter_i_14 ));
    CascadeMux I__5075 (
            .O(N__31526),
            .I(N__31523));
    InMux I__5074 (
            .O(N__31523),
            .I(N__31520));
    LocalMux I__5073 (
            .O(N__31520),
            .I(N__31517));
    Odrv12 I__5072 (
            .O(N__31517),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ));
    InMux I__5071 (
            .O(N__31514),
            .I(N__31511));
    LocalMux I__5070 (
            .O(N__31511),
            .I(\phase_controller_inst1.stoper_hc.counter_i_15 ));
    InMux I__5069 (
            .O(N__31508),
            .I(N__31505));
    LocalMux I__5068 (
            .O(N__31505),
            .I(N__31502));
    Odrv12 I__5067 (
            .O(N__31502),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ));
    CascadeMux I__5066 (
            .O(N__31499),
            .I(N__31496));
    InMux I__5065 (
            .O(N__31496),
            .I(N__31493));
    LocalMux I__5064 (
            .O(N__31493),
            .I(N__31490));
    Odrv12 I__5063 (
            .O(N__31490),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt20 ));
    CascadeMux I__5062 (
            .O(N__31487),
            .I(N__31484));
    InMux I__5061 (
            .O(N__31484),
            .I(N__31481));
    LocalMux I__5060 (
            .O(N__31481),
            .I(N__31478));
    Odrv4 I__5059 (
            .O(N__31478),
            .I(\phase_controller_inst1.stoper_hc.counter_i_3 ));
    CascadeMux I__5058 (
            .O(N__31475),
            .I(N__31472));
    InMux I__5057 (
            .O(N__31472),
            .I(N__31469));
    LocalMux I__5056 (
            .O(N__31469),
            .I(N__31466));
    Odrv4 I__5055 (
            .O(N__31466),
            .I(\phase_controller_inst1.stoper_hc.counter_i_4 ));
    InMux I__5054 (
            .O(N__31463),
            .I(N__31460));
    LocalMux I__5053 (
            .O(N__31460),
            .I(N__31457));
    Span4Mux_v I__5052 (
            .O(N__31457),
            .I(N__31454));
    Odrv4 I__5051 (
            .O(N__31454),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ));
    CascadeMux I__5050 (
            .O(N__31451),
            .I(N__31448));
    InMux I__5049 (
            .O(N__31448),
            .I(N__31445));
    LocalMux I__5048 (
            .O(N__31445),
            .I(N__31442));
    Odrv12 I__5047 (
            .O(N__31442),
            .I(\phase_controller_inst1.stoper_hc.counter_i_5 ));
    InMux I__5046 (
            .O(N__31439),
            .I(N__31436));
    LocalMux I__5045 (
            .O(N__31436),
            .I(\phase_controller_inst1.stoper_hc.counter_i_6 ));
    InMux I__5044 (
            .O(N__31433),
            .I(N__31430));
    LocalMux I__5043 (
            .O(N__31430),
            .I(\phase_controller_inst1.stoper_hc.counter_i_7 ));
    InMux I__5042 (
            .O(N__31427),
            .I(N__31424));
    LocalMux I__5041 (
            .O(N__31424),
            .I(N__31421));
    Odrv12 I__5040 (
            .O(N__31421),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ));
    CascadeMux I__5039 (
            .O(N__31418),
            .I(N__31415));
    InMux I__5038 (
            .O(N__31415),
            .I(N__31412));
    LocalMux I__5037 (
            .O(N__31412),
            .I(\phase_controller_inst1.stoper_hc.counter_i_8 ));
    InMux I__5036 (
            .O(N__31409),
            .I(N__31406));
    LocalMux I__5035 (
            .O(N__31406),
            .I(N__31403));
    Odrv12 I__5034 (
            .O(N__31403),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ));
    CascadeMux I__5033 (
            .O(N__31400),
            .I(N__31397));
    InMux I__5032 (
            .O(N__31397),
            .I(N__31394));
    LocalMux I__5031 (
            .O(N__31394),
            .I(\phase_controller_inst1.stoper_hc.counter_i_9 ));
    CascadeMux I__5030 (
            .O(N__31391),
            .I(N__31388));
    InMux I__5029 (
            .O(N__31388),
            .I(N__31385));
    LocalMux I__5028 (
            .O(N__31385),
            .I(\phase_controller_inst1.stoper_hc.counter_i_10 ));
    InMux I__5027 (
            .O(N__31382),
            .I(N__31376));
    InMux I__5026 (
            .O(N__31381),
            .I(N__31376));
    LocalMux I__5025 (
            .O(N__31376),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ));
    InMux I__5024 (
            .O(N__31373),
            .I(N__31367));
    InMux I__5023 (
            .O(N__31372),
            .I(N__31367));
    LocalMux I__5022 (
            .O(N__31367),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ));
    InMux I__5021 (
            .O(N__31364),
            .I(N__31358));
    InMux I__5020 (
            .O(N__31363),
            .I(N__31358));
    LocalMux I__5019 (
            .O(N__31358),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ));
    CascadeMux I__5018 (
            .O(N__31355),
            .I(N__31352));
    InMux I__5017 (
            .O(N__31352),
            .I(N__31349));
    LocalMux I__5016 (
            .O(N__31349),
            .I(\phase_controller_inst1.stoper_hc.counter_i_0 ));
    CascadeMux I__5015 (
            .O(N__31346),
            .I(N__31343));
    InMux I__5014 (
            .O(N__31343),
            .I(N__31340));
    LocalMux I__5013 (
            .O(N__31340),
            .I(N__31337));
    Span4Mux_v I__5012 (
            .O(N__31337),
            .I(N__31334));
    Odrv4 I__5011 (
            .O(N__31334),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ));
    InMux I__5010 (
            .O(N__31331),
            .I(N__31328));
    LocalMux I__5009 (
            .O(N__31328),
            .I(\phase_controller_inst1.stoper_hc.counter_i_1 ));
    CascadeMux I__5008 (
            .O(N__31325),
            .I(N__31322));
    InMux I__5007 (
            .O(N__31322),
            .I(N__31319));
    LocalMux I__5006 (
            .O(N__31319),
            .I(\phase_controller_inst1.stoper_hc.counter_i_2 ));
    InMux I__5005 (
            .O(N__31316),
            .I(N__31310));
    InMux I__5004 (
            .O(N__31315),
            .I(N__31310));
    LocalMux I__5003 (
            .O(N__31310),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ));
    InMux I__5002 (
            .O(N__31307),
            .I(N__31301));
    InMux I__5001 (
            .O(N__31306),
            .I(N__31301));
    LocalMux I__5000 (
            .O(N__31301),
            .I(N__31298));
    Odrv4 I__4999 (
            .O(N__31298),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ));
    InMux I__4998 (
            .O(N__31295),
            .I(N__31289));
    InMux I__4997 (
            .O(N__31294),
            .I(N__31289));
    LocalMux I__4996 (
            .O(N__31289),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ));
    InMux I__4995 (
            .O(N__31286),
            .I(N__31280));
    InMux I__4994 (
            .O(N__31285),
            .I(N__31280));
    LocalMux I__4993 (
            .O(N__31280),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ));
    InMux I__4992 (
            .O(N__31277),
            .I(N__31271));
    InMux I__4991 (
            .O(N__31276),
            .I(N__31271));
    LocalMux I__4990 (
            .O(N__31271),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ));
    InMux I__4989 (
            .O(N__31268),
            .I(N__31262));
    InMux I__4988 (
            .O(N__31267),
            .I(N__31262));
    LocalMux I__4987 (
            .O(N__31262),
            .I(N__31259));
    Odrv4 I__4986 (
            .O(N__31259),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ));
    InMux I__4985 (
            .O(N__31256),
            .I(N__31250));
    InMux I__4984 (
            .O(N__31255),
            .I(N__31250));
    LocalMux I__4983 (
            .O(N__31250),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ));
    InMux I__4982 (
            .O(N__31247),
            .I(N__31241));
    InMux I__4981 (
            .O(N__31246),
            .I(N__31241));
    LocalMux I__4980 (
            .O(N__31241),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ));
    InMux I__4979 (
            .O(N__31238),
            .I(N__31235));
    LocalMux I__4978 (
            .O(N__31235),
            .I(N__31231));
    InMux I__4977 (
            .O(N__31234),
            .I(N__31228));
    Span4Mux_h I__4976 (
            .O(N__31231),
            .I(N__31225));
    LocalMux I__4975 (
            .O(N__31228),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ));
    Odrv4 I__4974 (
            .O(N__31225),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ));
    InMux I__4973 (
            .O(N__31220),
            .I(N__31214));
    InMux I__4972 (
            .O(N__31219),
            .I(N__31214));
    LocalMux I__4971 (
            .O(N__31214),
            .I(N__31211));
    Odrv4 I__4970 (
            .O(N__31211),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ));
    CascadeMux I__4969 (
            .O(N__31208),
            .I(N__31204));
    CascadeMux I__4968 (
            .O(N__31207),
            .I(N__31201));
    InMux I__4967 (
            .O(N__31204),
            .I(N__31196));
    InMux I__4966 (
            .O(N__31201),
            .I(N__31196));
    LocalMux I__4965 (
            .O(N__31196),
            .I(N__31193));
    Odrv4 I__4964 (
            .O(N__31193),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ));
    CascadeMux I__4963 (
            .O(N__31190),
            .I(N__31186));
    CascadeMux I__4962 (
            .O(N__31189),
            .I(N__31183));
    InMux I__4961 (
            .O(N__31186),
            .I(N__31178));
    InMux I__4960 (
            .O(N__31183),
            .I(N__31178));
    LocalMux I__4959 (
            .O(N__31178),
            .I(N__31175));
    Odrv4 I__4958 (
            .O(N__31175),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ));
    InMux I__4957 (
            .O(N__31172),
            .I(N__31169));
    LocalMux I__4956 (
            .O(N__31169),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ));
    CascadeMux I__4955 (
            .O(N__31166),
            .I(N__31163));
    InMux I__4954 (
            .O(N__31163),
            .I(N__31160));
    LocalMux I__4953 (
            .O(N__31160),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt26 ));
    InMux I__4952 (
            .O(N__31157),
            .I(N__31154));
    LocalMux I__4951 (
            .O(N__31154),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt28 ));
    CascadeMux I__4950 (
            .O(N__31151),
            .I(N__31148));
    InMux I__4949 (
            .O(N__31148),
            .I(N__31145));
    LocalMux I__4948 (
            .O(N__31145),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ));
    InMux I__4947 (
            .O(N__31142),
            .I(N__31139));
    LocalMux I__4946 (
            .O(N__31139),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt30 ));
    CascadeMux I__4945 (
            .O(N__31136),
            .I(N__31133));
    InMux I__4944 (
            .O(N__31133),
            .I(N__31130));
    LocalMux I__4943 (
            .O(N__31130),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ));
    InMux I__4942 (
            .O(N__31127),
            .I(bfn_11_7_0_));
    CascadeMux I__4941 (
            .O(N__31124),
            .I(N__31119));
    InMux I__4940 (
            .O(N__31123),
            .I(N__31116));
    InMux I__4939 (
            .O(N__31122),
            .I(N__31111));
    InMux I__4938 (
            .O(N__31119),
            .I(N__31111));
    LocalMux I__4937 (
            .O(N__31116),
            .I(N__31108));
    LocalMux I__4936 (
            .O(N__31111),
            .I(N__31105));
    Span4Mux_s2_v I__4935 (
            .O(N__31108),
            .I(N__31102));
    Odrv4 I__4934 (
            .O(N__31105),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ));
    Odrv4 I__4933 (
            .O(N__31102),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ));
    InMux I__4932 (
            .O(N__31097),
            .I(N__31093));
    InMux I__4931 (
            .O(N__31096),
            .I(N__31090));
    LocalMux I__4930 (
            .O(N__31093),
            .I(N__31087));
    LocalMux I__4929 (
            .O(N__31090),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ));
    Odrv4 I__4928 (
            .O(N__31087),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ));
    CascadeMux I__4927 (
            .O(N__31082),
            .I(N__31079));
    InMux I__4926 (
            .O(N__31079),
            .I(N__31076));
    LocalMux I__4925 (
            .O(N__31076),
            .I(N__31073));
    Odrv4 I__4924 (
            .O(N__31073),
            .I(\phase_controller_inst2.stoper_hc.counter_i_13 ));
    InMux I__4923 (
            .O(N__31070),
            .I(N__31066));
    InMux I__4922 (
            .O(N__31069),
            .I(N__31063));
    LocalMux I__4921 (
            .O(N__31066),
            .I(N__31060));
    LocalMux I__4920 (
            .O(N__31063),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ));
    Odrv4 I__4919 (
            .O(N__31060),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ));
    CascadeMux I__4918 (
            .O(N__31055),
            .I(N__31052));
    InMux I__4917 (
            .O(N__31052),
            .I(N__31049));
    LocalMux I__4916 (
            .O(N__31049),
            .I(\phase_controller_inst2.stoper_hc.counter_i_14 ));
    InMux I__4915 (
            .O(N__31046),
            .I(N__31042));
    InMux I__4914 (
            .O(N__31045),
            .I(N__31039));
    LocalMux I__4913 (
            .O(N__31042),
            .I(N__31036));
    LocalMux I__4912 (
            .O(N__31039),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ));
    Odrv4 I__4911 (
            .O(N__31036),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ));
    InMux I__4910 (
            .O(N__31031),
            .I(N__31028));
    LocalMux I__4909 (
            .O(N__31028),
            .I(\phase_controller_inst2.stoper_hc.counter_i_15 ));
    InMux I__4908 (
            .O(N__31025),
            .I(N__31022));
    LocalMux I__4907 (
            .O(N__31022),
            .I(N__31019));
    Span4Mux_h I__4906 (
            .O(N__31019),
            .I(N__31016));
    Odrv4 I__4905 (
            .O(N__31016),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt16 ));
    CascadeMux I__4904 (
            .O(N__31013),
            .I(N__31010));
    InMux I__4903 (
            .O(N__31010),
            .I(N__31007));
    LocalMux I__4902 (
            .O(N__31007),
            .I(N__31004));
    Span4Mux_h I__4901 (
            .O(N__31004),
            .I(N__31001));
    Odrv4 I__4900 (
            .O(N__31001),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ));
    InMux I__4899 (
            .O(N__30998),
            .I(N__30995));
    LocalMux I__4898 (
            .O(N__30995),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ));
    CascadeMux I__4897 (
            .O(N__30992),
            .I(N__30989));
    InMux I__4896 (
            .O(N__30989),
            .I(N__30986));
    LocalMux I__4895 (
            .O(N__30986),
            .I(N__30983));
    Span4Mux_h I__4894 (
            .O(N__30983),
            .I(N__30980));
    Odrv4 I__4893 (
            .O(N__30980),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt18 ));
    InMux I__4892 (
            .O(N__30977),
            .I(N__30974));
    LocalMux I__4891 (
            .O(N__30974),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt20 ));
    CascadeMux I__4890 (
            .O(N__30971),
            .I(N__30968));
    InMux I__4889 (
            .O(N__30968),
            .I(N__30965));
    LocalMux I__4888 (
            .O(N__30965),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ));
    InMux I__4887 (
            .O(N__30962),
            .I(N__30959));
    LocalMux I__4886 (
            .O(N__30959),
            .I(N__30956));
    Odrv4 I__4885 (
            .O(N__30956),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ));
    CascadeMux I__4884 (
            .O(N__30953),
            .I(N__30950));
    InMux I__4883 (
            .O(N__30950),
            .I(N__30947));
    LocalMux I__4882 (
            .O(N__30947),
            .I(N__30944));
    Odrv4 I__4881 (
            .O(N__30944),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt22 ));
    InMux I__4880 (
            .O(N__30941),
            .I(N__30938));
    LocalMux I__4879 (
            .O(N__30938),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ));
    CascadeMux I__4878 (
            .O(N__30935),
            .I(N__30932));
    InMux I__4877 (
            .O(N__30932),
            .I(N__30929));
    LocalMux I__4876 (
            .O(N__30929),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt24 ));
    InMux I__4875 (
            .O(N__30926),
            .I(N__30922));
    InMux I__4874 (
            .O(N__30925),
            .I(N__30919));
    LocalMux I__4873 (
            .O(N__30922),
            .I(N__30916));
    LocalMux I__4872 (
            .O(N__30919),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ));
    Odrv4 I__4871 (
            .O(N__30916),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ));
    InMux I__4870 (
            .O(N__30911),
            .I(N__30908));
    LocalMux I__4869 (
            .O(N__30908),
            .I(\phase_controller_inst2.stoper_hc.counter_i_5 ));
    InMux I__4868 (
            .O(N__30905),
            .I(N__30901));
    InMux I__4867 (
            .O(N__30904),
            .I(N__30898));
    LocalMux I__4866 (
            .O(N__30901),
            .I(N__30895));
    LocalMux I__4865 (
            .O(N__30898),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ));
    Odrv4 I__4864 (
            .O(N__30895),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ));
    InMux I__4863 (
            .O(N__30890),
            .I(N__30887));
    LocalMux I__4862 (
            .O(N__30887),
            .I(\phase_controller_inst2.stoper_hc.counter_i_6 ));
    InMux I__4861 (
            .O(N__30884),
            .I(N__30880));
    InMux I__4860 (
            .O(N__30883),
            .I(N__30877));
    LocalMux I__4859 (
            .O(N__30880),
            .I(N__30874));
    LocalMux I__4858 (
            .O(N__30877),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ));
    Odrv4 I__4857 (
            .O(N__30874),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ));
    InMux I__4856 (
            .O(N__30869),
            .I(N__30866));
    LocalMux I__4855 (
            .O(N__30866),
            .I(\phase_controller_inst2.stoper_hc.counter_i_7 ));
    InMux I__4854 (
            .O(N__30863),
            .I(N__30860));
    LocalMux I__4853 (
            .O(N__30860),
            .I(N__30856));
    InMux I__4852 (
            .O(N__30859),
            .I(N__30853));
    Span4Mux_v I__4851 (
            .O(N__30856),
            .I(N__30850));
    LocalMux I__4850 (
            .O(N__30853),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ));
    Odrv4 I__4849 (
            .O(N__30850),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ));
    CascadeMux I__4848 (
            .O(N__30845),
            .I(N__30842));
    InMux I__4847 (
            .O(N__30842),
            .I(N__30839));
    LocalMux I__4846 (
            .O(N__30839),
            .I(\phase_controller_inst2.stoper_hc.counter_i_8 ));
    InMux I__4845 (
            .O(N__30836),
            .I(N__30832));
    InMux I__4844 (
            .O(N__30835),
            .I(N__30829));
    LocalMux I__4843 (
            .O(N__30832),
            .I(N__30826));
    LocalMux I__4842 (
            .O(N__30829),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ));
    Odrv4 I__4841 (
            .O(N__30826),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ));
    InMux I__4840 (
            .O(N__30821),
            .I(N__30818));
    LocalMux I__4839 (
            .O(N__30818),
            .I(\phase_controller_inst2.stoper_hc.counter_i_9 ));
    InMux I__4838 (
            .O(N__30815),
            .I(N__30812));
    LocalMux I__4837 (
            .O(N__30812),
            .I(N__30808));
    InMux I__4836 (
            .O(N__30811),
            .I(N__30805));
    Span4Mux_v I__4835 (
            .O(N__30808),
            .I(N__30802));
    LocalMux I__4834 (
            .O(N__30805),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ));
    Odrv4 I__4833 (
            .O(N__30802),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ));
    CascadeMux I__4832 (
            .O(N__30797),
            .I(N__30794));
    InMux I__4831 (
            .O(N__30794),
            .I(N__30791));
    LocalMux I__4830 (
            .O(N__30791),
            .I(\phase_controller_inst2.stoper_hc.counter_i_10 ));
    InMux I__4829 (
            .O(N__30788),
            .I(N__30784));
    InMux I__4828 (
            .O(N__30787),
            .I(N__30781));
    LocalMux I__4827 (
            .O(N__30784),
            .I(N__30778));
    LocalMux I__4826 (
            .O(N__30781),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ));
    Odrv4 I__4825 (
            .O(N__30778),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ));
    CascadeMux I__4824 (
            .O(N__30773),
            .I(N__30770));
    InMux I__4823 (
            .O(N__30770),
            .I(N__30767));
    LocalMux I__4822 (
            .O(N__30767),
            .I(N__30764));
    Odrv4 I__4821 (
            .O(N__30764),
            .I(\phase_controller_inst2.stoper_hc.counter_i_11 ));
    InMux I__4820 (
            .O(N__30761),
            .I(N__30757));
    InMux I__4819 (
            .O(N__30760),
            .I(N__30754));
    LocalMux I__4818 (
            .O(N__30757),
            .I(N__30751));
    LocalMux I__4817 (
            .O(N__30754),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ));
    Odrv4 I__4816 (
            .O(N__30751),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ));
    CascadeMux I__4815 (
            .O(N__30746),
            .I(N__30743));
    InMux I__4814 (
            .O(N__30743),
            .I(N__30740));
    LocalMux I__4813 (
            .O(N__30740),
            .I(\phase_controller_inst2.stoper_hc.counter_i_12 ));
    InMux I__4812 (
            .O(N__30737),
            .I(N__30734));
    LocalMux I__4811 (
            .O(N__30734),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    CascadeMux I__4810 (
            .O(N__30731),
            .I(N__30726));
    InMux I__4809 (
            .O(N__30730),
            .I(N__30723));
    InMux I__4808 (
            .O(N__30729),
            .I(N__30717));
    InMux I__4807 (
            .O(N__30726),
            .I(N__30717));
    LocalMux I__4806 (
            .O(N__30723),
            .I(N__30714));
    InMux I__4805 (
            .O(N__30722),
            .I(N__30711));
    LocalMux I__4804 (
            .O(N__30717),
            .I(N__30708));
    Span12Mux_s11_v I__4803 (
            .O(N__30714),
            .I(N__30705));
    LocalMux I__4802 (
            .O(N__30711),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__4801 (
            .O(N__30708),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__4800 (
            .O(N__30705),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__4799 (
            .O(N__30698),
            .I(N__30695));
    LocalMux I__4798 (
            .O(N__30695),
            .I(N__30692));
    Span4Mux_s2_v I__4797 (
            .O(N__30692),
            .I(N__30689));
    Odrv4 I__4796 (
            .O(N__30689),
            .I(s2_phy_c));
    InMux I__4795 (
            .O(N__30686),
            .I(N__30679));
    CascadeMux I__4794 (
            .O(N__30685),
            .I(N__30676));
    InMux I__4793 (
            .O(N__30684),
            .I(N__30672));
    InMux I__4792 (
            .O(N__30683),
            .I(N__30667));
    InMux I__4791 (
            .O(N__30682),
            .I(N__30667));
    LocalMux I__4790 (
            .O(N__30679),
            .I(N__30664));
    InMux I__4789 (
            .O(N__30676),
            .I(N__30661));
    InMux I__4788 (
            .O(N__30675),
            .I(N__30658));
    LocalMux I__4787 (
            .O(N__30672),
            .I(N__30655));
    LocalMux I__4786 (
            .O(N__30667),
            .I(N__30652));
    Span12Mux_s6_v I__4785 (
            .O(N__30664),
            .I(N__30649));
    LocalMux I__4784 (
            .O(N__30661),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__4783 (
            .O(N__30658),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv12 I__4782 (
            .O(N__30655),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__4781 (
            .O(N__30652),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv12 I__4780 (
            .O(N__30649),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    CascadeMux I__4779 (
            .O(N__30638),
            .I(N__30634));
    InMux I__4778 (
            .O(N__30637),
            .I(N__30631));
    InMux I__4777 (
            .O(N__30634),
            .I(N__30628));
    LocalMux I__4776 (
            .O(N__30631),
            .I(\phase_controller_inst2.stoper_hc.counter ));
    LocalMux I__4775 (
            .O(N__30628),
            .I(\phase_controller_inst2.stoper_hc.counter ));
    InMux I__4774 (
            .O(N__30623),
            .I(N__30620));
    LocalMux I__4773 (
            .O(N__30620),
            .I(N__30616));
    InMux I__4772 (
            .O(N__30619),
            .I(N__30613));
    Span4Mux_v I__4771 (
            .O(N__30616),
            .I(N__30610));
    LocalMux I__4770 (
            .O(N__30613),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ));
    Odrv4 I__4769 (
            .O(N__30610),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ));
    InMux I__4768 (
            .O(N__30605),
            .I(N__30602));
    LocalMux I__4767 (
            .O(N__30602),
            .I(\phase_controller_inst2.stoper_hc.counter_i_0 ));
    InMux I__4766 (
            .O(N__30599),
            .I(N__30595));
    InMux I__4765 (
            .O(N__30598),
            .I(N__30592));
    LocalMux I__4764 (
            .O(N__30595),
            .I(N__30589));
    LocalMux I__4763 (
            .O(N__30592),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ));
    Odrv4 I__4762 (
            .O(N__30589),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ));
    CascadeMux I__4761 (
            .O(N__30584),
            .I(N__30581));
    InMux I__4760 (
            .O(N__30581),
            .I(N__30578));
    LocalMux I__4759 (
            .O(N__30578),
            .I(\phase_controller_inst2.stoper_hc.counter_i_1 ));
    InMux I__4758 (
            .O(N__30575),
            .I(N__30572));
    LocalMux I__4757 (
            .O(N__30572),
            .I(N__30568));
    InMux I__4756 (
            .O(N__30571),
            .I(N__30565));
    Span4Mux_v I__4755 (
            .O(N__30568),
            .I(N__30562));
    LocalMux I__4754 (
            .O(N__30565),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ));
    Odrv4 I__4753 (
            .O(N__30562),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ));
    CascadeMux I__4752 (
            .O(N__30557),
            .I(N__30554));
    InMux I__4751 (
            .O(N__30554),
            .I(N__30551));
    LocalMux I__4750 (
            .O(N__30551),
            .I(\phase_controller_inst2.stoper_hc.counter_i_2 ));
    InMux I__4749 (
            .O(N__30548),
            .I(N__30544));
    InMux I__4748 (
            .O(N__30547),
            .I(N__30541));
    LocalMux I__4747 (
            .O(N__30544),
            .I(N__30538));
    LocalMux I__4746 (
            .O(N__30541),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ));
    Odrv4 I__4745 (
            .O(N__30538),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ));
    InMux I__4744 (
            .O(N__30533),
            .I(N__30530));
    LocalMux I__4743 (
            .O(N__30530),
            .I(\phase_controller_inst2.stoper_hc.counter_i_3 ));
    InMux I__4742 (
            .O(N__30527),
            .I(N__30523));
    InMux I__4741 (
            .O(N__30526),
            .I(N__30520));
    LocalMux I__4740 (
            .O(N__30523),
            .I(N__30517));
    LocalMux I__4739 (
            .O(N__30520),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ));
    Odrv4 I__4738 (
            .O(N__30517),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ));
    CascadeMux I__4737 (
            .O(N__30512),
            .I(N__30509));
    InMux I__4736 (
            .O(N__30509),
            .I(N__30506));
    LocalMux I__4735 (
            .O(N__30506),
            .I(\phase_controller_inst2.stoper_hc.counter_i_4 ));
    InMux I__4734 (
            .O(N__30503),
            .I(N__30500));
    LocalMux I__4733 (
            .O(N__30500),
            .I(N__30496));
    InMux I__4732 (
            .O(N__30499),
            .I(N__30493));
    Odrv4 I__4731 (
            .O(N__30496),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ));
    LocalMux I__4730 (
            .O(N__30493),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ));
    InMux I__4729 (
            .O(N__30488),
            .I(N__30484));
    InMux I__4728 (
            .O(N__30487),
            .I(N__30481));
    LocalMux I__4727 (
            .O(N__30484),
            .I(N__30477));
    LocalMux I__4726 (
            .O(N__30481),
            .I(N__30474));
    InMux I__4725 (
            .O(N__30480),
            .I(N__30471));
    Span4Mux_v I__4724 (
            .O(N__30477),
            .I(N__30466));
    Span4Mux_v I__4723 (
            .O(N__30474),
            .I(N__30466));
    LocalMux I__4722 (
            .O(N__30471),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ));
    Odrv4 I__4721 (
            .O(N__30466),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ));
    CascadeMux I__4720 (
            .O(N__30461),
            .I(N__30458));
    InMux I__4719 (
            .O(N__30458),
            .I(N__30454));
    InMux I__4718 (
            .O(N__30457),
            .I(N__30451));
    LocalMux I__4717 (
            .O(N__30454),
            .I(N__30448));
    LocalMux I__4716 (
            .O(N__30451),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ));
    Odrv4 I__4715 (
            .O(N__30448),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ));
    CascadeMux I__4714 (
            .O(N__30443),
            .I(N__30439));
    InMux I__4713 (
            .O(N__30442),
            .I(N__30436));
    InMux I__4712 (
            .O(N__30439),
            .I(N__30433));
    LocalMux I__4711 (
            .O(N__30436),
            .I(N__30427));
    LocalMux I__4710 (
            .O(N__30433),
            .I(N__30427));
    InMux I__4709 (
            .O(N__30432),
            .I(N__30424));
    Span4Mux_v I__4708 (
            .O(N__30427),
            .I(N__30421));
    LocalMux I__4707 (
            .O(N__30424),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ));
    Odrv4 I__4706 (
            .O(N__30421),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ));
    InMux I__4705 (
            .O(N__30416),
            .I(N__30413));
    LocalMux I__4704 (
            .O(N__30413),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt20 ));
    InMux I__4703 (
            .O(N__30410),
            .I(N__30407));
    LocalMux I__4702 (
            .O(N__30407),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    CascadeMux I__4701 (
            .O(N__30404),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_));
    InMux I__4700 (
            .O(N__30401),
            .I(N__30398));
    LocalMux I__4699 (
            .O(N__30398),
            .I(N__30395));
    Span4Mux_h I__4698 (
            .O(N__30395),
            .I(N__30392));
    Span4Mux_v I__4697 (
            .O(N__30392),
            .I(N__30389));
    Odrv4 I__4696 (
            .O(N__30389),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ));
    InMux I__4695 (
            .O(N__30386),
            .I(N__30382));
    InMux I__4694 (
            .O(N__30385),
            .I(N__30379));
    LocalMux I__4693 (
            .O(N__30382),
            .I(N__30374));
    LocalMux I__4692 (
            .O(N__30379),
            .I(N__30374));
    Odrv4 I__4691 (
            .O(N__30374),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ));
    InMux I__4690 (
            .O(N__30371),
            .I(N__30368));
    LocalMux I__4689 (
            .O(N__30368),
            .I(N__30364));
    InMux I__4688 (
            .O(N__30367),
            .I(N__30360));
    Span4Mux_h I__4687 (
            .O(N__30364),
            .I(N__30357));
    InMux I__4686 (
            .O(N__30363),
            .I(N__30354));
    LocalMux I__4685 (
            .O(N__30360),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ));
    Odrv4 I__4684 (
            .O(N__30357),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ));
    LocalMux I__4683 (
            .O(N__30354),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ));
    CascadeMux I__4682 (
            .O(N__30347),
            .I(N__30344));
    InMux I__4681 (
            .O(N__30344),
            .I(N__30340));
    CascadeMux I__4680 (
            .O(N__30343),
            .I(N__30336));
    LocalMux I__4679 (
            .O(N__30340),
            .I(N__30333));
    InMux I__4678 (
            .O(N__30339),
            .I(N__30330));
    InMux I__4677 (
            .O(N__30336),
            .I(N__30327));
    Span4Mux_h I__4676 (
            .O(N__30333),
            .I(N__30324));
    LocalMux I__4675 (
            .O(N__30330),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ));
    LocalMux I__4674 (
            .O(N__30327),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ));
    Odrv4 I__4673 (
            .O(N__30324),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ));
    InMux I__4672 (
            .O(N__30317),
            .I(N__30313));
    InMux I__4671 (
            .O(N__30316),
            .I(N__30310));
    LocalMux I__4670 (
            .O(N__30313),
            .I(N__30305));
    LocalMux I__4669 (
            .O(N__30310),
            .I(N__30305));
    Odrv4 I__4668 (
            .O(N__30305),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ));
    CascadeMux I__4667 (
            .O(N__30302),
            .I(N__30299));
    InMux I__4666 (
            .O(N__30299),
            .I(N__30296));
    LocalMux I__4665 (
            .O(N__30296),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt22 ));
    InMux I__4664 (
            .O(N__30293),
            .I(N__30290));
    LocalMux I__4663 (
            .O(N__30290),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    CascadeMux I__4662 (
            .O(N__30287),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ));
    InMux I__4661 (
            .O(N__30284),
            .I(N__30281));
    LocalMux I__4660 (
            .O(N__30281),
            .I(N__30278));
    Span12Mux_v I__4659 (
            .O(N__30278),
            .I(N__30275));
    Odrv12 I__4658 (
            .O(N__30275),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    InMux I__4657 (
            .O(N__30272),
            .I(N__30269));
    LocalMux I__4656 (
            .O(N__30269),
            .I(N__30266));
    Span4Mux_h I__4655 (
            .O(N__30266),
            .I(N__30263));
    Sp12to4 I__4654 (
            .O(N__30263),
            .I(N__30260));
    Span12Mux_v I__4653 (
            .O(N__30260),
            .I(N__30257));
    Odrv12 I__4652 (
            .O(N__30257),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__4651 (
            .O(N__30254),
            .I(N__30251));
    LocalMux I__4650 (
            .O(N__30251),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    CascadeMux I__4649 (
            .O(N__30248),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_));
    InMux I__4648 (
            .O(N__30245),
            .I(N__30242));
    LocalMux I__4647 (
            .O(N__30242),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ));
    InMux I__4646 (
            .O(N__30239),
            .I(N__30235));
    InMux I__4645 (
            .O(N__30238),
            .I(N__30232));
    LocalMux I__4644 (
            .O(N__30235),
            .I(N__30229));
    LocalMux I__4643 (
            .O(N__30232),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_20));
    Odrv4 I__4642 (
            .O(N__30229),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_20));
    InMux I__4641 (
            .O(N__30224),
            .I(N__30220));
    InMux I__4640 (
            .O(N__30223),
            .I(N__30217));
    LocalMux I__4639 (
            .O(N__30220),
            .I(N__30214));
    LocalMux I__4638 (
            .O(N__30217),
            .I(N__30211));
    Odrv4 I__4637 (
            .O(N__30214),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_21));
    Odrv4 I__4636 (
            .O(N__30211),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_21));
    InMux I__4635 (
            .O(N__30206),
            .I(N__30202));
    InMux I__4634 (
            .O(N__30205),
            .I(N__30199));
    LocalMux I__4633 (
            .O(N__30202),
            .I(N__30196));
    LocalMux I__4632 (
            .O(N__30199),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_22));
    Odrv4 I__4631 (
            .O(N__30196),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_22));
    InMux I__4630 (
            .O(N__30191),
            .I(N__30188));
    LocalMux I__4629 (
            .O(N__30188),
            .I(N__30185));
    Span4Mux_v I__4628 (
            .O(N__30185),
            .I(N__30181));
    InMux I__4627 (
            .O(N__30184),
            .I(N__30178));
    Span4Mux_v I__4626 (
            .O(N__30181),
            .I(N__30173));
    LocalMux I__4625 (
            .O(N__30178),
            .I(N__30173));
    Odrv4 I__4624 (
            .O(N__30173),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_23));
    CascadeMux I__4623 (
            .O(N__30170),
            .I(N__30167));
    InMux I__4622 (
            .O(N__30167),
            .I(N__30164));
    LocalMux I__4621 (
            .O(N__30164),
            .I(N__30161));
    Odrv4 I__4620 (
            .O(N__30161),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ));
    InMux I__4619 (
            .O(N__30158),
            .I(N__30155));
    LocalMux I__4618 (
            .O(N__30155),
            .I(N__30152));
    Span4Mux_v I__4617 (
            .O(N__30152),
            .I(N__30149));
    Odrv4 I__4616 (
            .O(N__30149),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ));
    CascadeMux I__4615 (
            .O(N__30146),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ));
    InMux I__4614 (
            .O(N__30143),
            .I(N__30140));
    LocalMux I__4613 (
            .O(N__30140),
            .I(N__30137));
    Odrv12 I__4612 (
            .O(N__30137),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ));
    InMux I__4611 (
            .O(N__30134),
            .I(N__30131));
    LocalMux I__4610 (
            .O(N__30131),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ));
    InMux I__4609 (
            .O(N__30128),
            .I(N__30125));
    LocalMux I__4608 (
            .O(N__30125),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    CascadeMux I__4607 (
            .O(N__30122),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_));
    InMux I__4606 (
            .O(N__30119),
            .I(N__30116));
    LocalMux I__4605 (
            .O(N__30116),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ));
    InMux I__4604 (
            .O(N__30113),
            .I(N__30109));
    InMux I__4603 (
            .O(N__30112),
            .I(N__30106));
    LocalMux I__4602 (
            .O(N__30109),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    LocalMux I__4601 (
            .O(N__30106),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__4600 (
            .O(N__30101),
            .I(N__30098));
    LocalMux I__4599 (
            .O(N__30098),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    CascadeMux I__4598 (
            .O(N__30095),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_));
    InMux I__4597 (
            .O(N__30092),
            .I(N__30089));
    LocalMux I__4596 (
            .O(N__30089),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ));
    InMux I__4595 (
            .O(N__30086),
            .I(N__30083));
    LocalMux I__4594 (
            .O(N__30083),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    CascadeMux I__4593 (
            .O(N__30080),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_));
    InMux I__4592 (
            .O(N__30077),
            .I(N__30074));
    LocalMux I__4591 (
            .O(N__30074),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ));
    InMux I__4590 (
            .O(N__30071),
            .I(N__30068));
    LocalMux I__4589 (
            .O(N__30068),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    CascadeMux I__4588 (
            .O(N__30065),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_));
    InMux I__4587 (
            .O(N__30062),
            .I(N__30059));
    LocalMux I__4586 (
            .O(N__30059),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ));
    InMux I__4585 (
            .O(N__30056),
            .I(N__30052));
    InMux I__4584 (
            .O(N__30055),
            .I(N__30049));
    LocalMux I__4583 (
            .O(N__30052),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__4582 (
            .O(N__30049),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    InMux I__4581 (
            .O(N__30044),
            .I(N__30041));
    LocalMux I__4580 (
            .O(N__30041),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ));
    InMux I__4579 (
            .O(N__30038),
            .I(N__30035));
    LocalMux I__4578 (
            .O(N__30035),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    CascadeMux I__4577 (
            .O(N__30032),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_));
    InMux I__4576 (
            .O(N__30029),
            .I(N__30026));
    LocalMux I__4575 (
            .O(N__30026),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ));
    InMux I__4574 (
            .O(N__30023),
            .I(N__30020));
    LocalMux I__4573 (
            .O(N__30020),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    CascadeMux I__4572 (
            .O(N__30017),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17_cascade_));
    CascadeMux I__4571 (
            .O(N__30014),
            .I(N__30011));
    InMux I__4570 (
            .O(N__30011),
            .I(N__30008));
    LocalMux I__4569 (
            .O(N__30008),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ));
    InMux I__4568 (
            .O(N__30005),
            .I(N__30001));
    InMux I__4567 (
            .O(N__30004),
            .I(N__29998));
    LocalMux I__4566 (
            .O(N__30001),
            .I(N__29995));
    LocalMux I__4565 (
            .O(N__29998),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    Odrv12 I__4564 (
            .O(N__29995),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    InMux I__4563 (
            .O(N__29990),
            .I(N__29987));
    LocalMux I__4562 (
            .O(N__29987),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ));
    InMux I__4561 (
            .O(N__29984),
            .I(N__29981));
    LocalMux I__4560 (
            .O(N__29981),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    CascadeMux I__4559 (
            .O(N__29978),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_));
    InMux I__4558 (
            .O(N__29975),
            .I(N__29972));
    LocalMux I__4557 (
            .O(N__29972),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    CascadeMux I__4556 (
            .O(N__29969),
            .I(elapsed_time_ns_1_RNIGF91B_0_4_cascade_));
    InMux I__4555 (
            .O(N__29966),
            .I(N__29963));
    LocalMux I__4554 (
            .O(N__29963),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ));
    InMux I__4553 (
            .O(N__29960),
            .I(N__29956));
    InMux I__4552 (
            .O(N__29959),
            .I(N__29953));
    LocalMux I__4551 (
            .O(N__29956),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__4550 (
            .O(N__29953),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    InMux I__4549 (
            .O(N__29948),
            .I(N__29945));
    LocalMux I__4548 (
            .O(N__29945),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ));
    InMux I__4547 (
            .O(N__29942),
            .I(N__29939));
    LocalMux I__4546 (
            .O(N__29939),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    CascadeMux I__4545 (
            .O(N__29936),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_));
    CascadeMux I__4544 (
            .O(N__29933),
            .I(N__29930));
    InMux I__4543 (
            .O(N__29930),
            .I(N__29927));
    LocalMux I__4542 (
            .O(N__29927),
            .I(N__29924));
    Odrv4 I__4541 (
            .O(N__29924),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ));
    InMux I__4540 (
            .O(N__29921),
            .I(N__29917));
    InMux I__4539 (
            .O(N__29920),
            .I(N__29914));
    LocalMux I__4538 (
            .O(N__29917),
            .I(N__29911));
    LocalMux I__4537 (
            .O(N__29914),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    Odrv4 I__4536 (
            .O(N__29911),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__4535 (
            .O(N__29906),
            .I(N__29903));
    LocalMux I__4534 (
            .O(N__29903),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ));
    InMux I__4533 (
            .O(N__29900),
            .I(N__29897));
    LocalMux I__4532 (
            .O(N__29897),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    CascadeMux I__4531 (
            .O(N__29894),
            .I(elapsed_time_ns_1_RNIHG91B_0_5_cascade_));
    InMux I__4530 (
            .O(N__29891),
            .I(N__29888));
    LocalMux I__4529 (
            .O(N__29888),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ));
    InMux I__4528 (
            .O(N__29885),
            .I(N__29882));
    LocalMux I__4527 (
            .O(N__29882),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__4526 (
            .O(N__29879),
            .I(N__29875));
    InMux I__4525 (
            .O(N__29878),
            .I(N__29872));
    LocalMux I__4524 (
            .O(N__29875),
            .I(N__29869));
    LocalMux I__4523 (
            .O(N__29872),
            .I(N__29866));
    Span12Mux_v I__4522 (
            .O(N__29869),
            .I(N__29863));
    Span12Mux_v I__4521 (
            .O(N__29866),
            .I(N__29860));
    Span12Mux_h I__4520 (
            .O(N__29863),
            .I(N__29857));
    Span12Mux_h I__4519 (
            .O(N__29860),
            .I(N__29854));
    Span12Mux_h I__4518 (
            .O(N__29857),
            .I(N__29851));
    Odrv12 I__4517 (
            .O(N__29854),
            .I(\pwm_generator_inst.un3_threshold ));
    Odrv12 I__4516 (
            .O(N__29851),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__4515 (
            .O(N__29846),
            .I(N__29843));
    LocalMux I__4514 (
            .O(N__29843),
            .I(N__29840));
    Span4Mux_h I__4513 (
            .O(N__29840),
            .I(N__29837));
    Sp12to4 I__4512 (
            .O(N__29837),
            .I(N__29834));
    Span12Mux_v I__4511 (
            .O(N__29834),
            .I(N__29831));
    Odrv12 I__4510 (
            .O(N__29831),
            .I(\pwm_generator_inst.un3_threshold_iZ0 ));
    InMux I__4509 (
            .O(N__29828),
            .I(N__29825));
    LocalMux I__4508 (
            .O(N__29825),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ));
    CascadeMux I__4507 (
            .O(N__29822),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ));
    CascadeMux I__4506 (
            .O(N__29819),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__4505 (
            .O(N__29816),
            .I(N__29813));
    LocalMux I__4504 (
            .O(N__29813),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    CascadeMux I__4503 (
            .O(N__29810),
            .I(elapsed_time_ns_1_RNIIH91B_0_6_cascade_));
    InMux I__4502 (
            .O(N__29807),
            .I(N__29804));
    LocalMux I__4501 (
            .O(N__29804),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ));
    InMux I__4500 (
            .O(N__29801),
            .I(N__29798));
    LocalMux I__4499 (
            .O(N__29798),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    CascadeMux I__4498 (
            .O(N__29795),
            .I(elapsed_time_ns_1_RNILK91B_0_9_cascade_));
    InMux I__4497 (
            .O(N__29792),
            .I(N__29789));
    LocalMux I__4496 (
            .O(N__29789),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ));
    InMux I__4495 (
            .O(N__29786),
            .I(N__29782));
    InMux I__4494 (
            .O(N__29785),
            .I(N__29779));
    LocalMux I__4493 (
            .O(N__29782),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    LocalMux I__4492 (
            .O(N__29779),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    InMux I__4491 (
            .O(N__29774),
            .I(N__29764));
    InMux I__4490 (
            .O(N__29773),
            .I(N__29764));
    InMux I__4489 (
            .O(N__29772),
            .I(N__29764));
    InMux I__4488 (
            .O(N__29771),
            .I(N__29761));
    LocalMux I__4487 (
            .O(N__29764),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__4486 (
            .O(N__29761),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__4485 (
            .O(N__29756),
            .I(N__29753));
    LocalMux I__4484 (
            .O(N__29753),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__4483 (
            .O(N__29750),
            .I(N__29747));
    LocalMux I__4482 (
            .O(N__29747),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    CascadeMux I__4481 (
            .O(N__29744),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_));
    InMux I__4480 (
            .O(N__29741),
            .I(N__29738));
    LocalMux I__4479 (
            .O(N__29738),
            .I(N__29735));
    Odrv4 I__4478 (
            .O(N__29735),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ));
    InMux I__4477 (
            .O(N__29732),
            .I(N__29729));
    LocalMux I__4476 (
            .O(N__29729),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    CascadeMux I__4475 (
            .O(N__29726),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8_cascade_));
    InMux I__4474 (
            .O(N__29723),
            .I(N__29720));
    LocalMux I__4473 (
            .O(N__29720),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ));
    InMux I__4472 (
            .O(N__29717),
            .I(N__29710));
    InMux I__4471 (
            .O(N__29716),
            .I(N__29710));
    InMux I__4470 (
            .O(N__29715),
            .I(N__29707));
    LocalMux I__4469 (
            .O(N__29710),
            .I(N__29704));
    LocalMux I__4468 (
            .O(N__29707),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ));
    Odrv12 I__4467 (
            .O(N__29704),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ));
    InMux I__4466 (
            .O(N__29699),
            .I(N__29693));
    InMux I__4465 (
            .O(N__29698),
            .I(N__29693));
    LocalMux I__4464 (
            .O(N__29693),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ));
    CascadeMux I__4463 (
            .O(N__29690),
            .I(N__29686));
    CascadeMux I__4462 (
            .O(N__29689),
            .I(N__29683));
    InMux I__4461 (
            .O(N__29686),
            .I(N__29677));
    InMux I__4460 (
            .O(N__29683),
            .I(N__29677));
    InMux I__4459 (
            .O(N__29682),
            .I(N__29674));
    LocalMux I__4458 (
            .O(N__29677),
            .I(N__29671));
    LocalMux I__4457 (
            .O(N__29674),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_16 ));
    Odrv12 I__4456 (
            .O(N__29671),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_16 ));
    InMux I__4455 (
            .O(N__29666),
            .I(N__29662));
    InMux I__4454 (
            .O(N__29665),
            .I(N__29659));
    LocalMux I__4453 (
            .O(N__29662),
            .I(N__29656));
    LocalMux I__4452 (
            .O(N__29659),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ));
    Odrv4 I__4451 (
            .O(N__29656),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ));
    InMux I__4450 (
            .O(N__29651),
            .I(N__29639));
    InMux I__4449 (
            .O(N__29650),
            .I(N__29639));
    InMux I__4448 (
            .O(N__29649),
            .I(N__29639));
    InMux I__4447 (
            .O(N__29648),
            .I(N__29639));
    LocalMux I__4446 (
            .O(N__29639),
            .I(N__29636));
    Span4Mux_h I__4445 (
            .O(N__29636),
            .I(N__29633));
    Odrv4 I__4444 (
            .O(N__29633),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ));
    InMux I__4443 (
            .O(N__29630),
            .I(N__29624));
    InMux I__4442 (
            .O(N__29629),
            .I(N__29624));
    LocalMux I__4441 (
            .O(N__29624),
            .I(N__29621));
    Odrv12 I__4440 (
            .O(N__29621),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ));
    InMux I__4439 (
            .O(N__29618),
            .I(N__29615));
    LocalMux I__4438 (
            .O(N__29615),
            .I(N__29610));
    InMux I__4437 (
            .O(N__29614),
            .I(N__29607));
    InMux I__4436 (
            .O(N__29613),
            .I(N__29604));
    Span12Mux_h I__4435 (
            .O(N__29610),
            .I(N__29597));
    LocalMux I__4434 (
            .O(N__29607),
            .I(N__29597));
    LocalMux I__4433 (
            .O(N__29604),
            .I(N__29597));
    Odrv12 I__4432 (
            .O(N__29597),
            .I(il_min_comp1_c));
    InMux I__4431 (
            .O(N__29594),
            .I(N__29587));
    InMux I__4430 (
            .O(N__29593),
            .I(N__29587));
    InMux I__4429 (
            .O(N__29592),
            .I(N__29584));
    LocalMux I__4428 (
            .O(N__29587),
            .I(N__29579));
    LocalMux I__4427 (
            .O(N__29584),
            .I(N__29579));
    Span4Mux_h I__4426 (
            .O(N__29579),
            .I(N__29576));
    Span4Mux_v I__4425 (
            .O(N__29576),
            .I(N__29573));
    Span4Mux_v I__4424 (
            .O(N__29573),
            .I(N__29570));
    Odrv4 I__4423 (
            .O(N__29570),
            .I(il_max_comp1_c));
    InMux I__4422 (
            .O(N__29567),
            .I(N__29560));
    InMux I__4421 (
            .O(N__29566),
            .I(N__29560));
    InMux I__4420 (
            .O(N__29565),
            .I(N__29557));
    LocalMux I__4419 (
            .O(N__29560),
            .I(N__29554));
    LocalMux I__4418 (
            .O(N__29557),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ));
    Odrv4 I__4417 (
            .O(N__29554),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ));
    InMux I__4416 (
            .O(N__29549),
            .I(N__29542));
    InMux I__4415 (
            .O(N__29548),
            .I(N__29542));
    InMux I__4414 (
            .O(N__29547),
            .I(N__29539));
    LocalMux I__4413 (
            .O(N__29542),
            .I(N__29536));
    LocalMux I__4412 (
            .O(N__29539),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ));
    Odrv4 I__4411 (
            .O(N__29536),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ));
    InMux I__4410 (
            .O(N__29531),
            .I(N__29524));
    InMux I__4409 (
            .O(N__29530),
            .I(N__29524));
    InMux I__4408 (
            .O(N__29529),
            .I(N__29521));
    LocalMux I__4407 (
            .O(N__29524),
            .I(N__29518));
    LocalMux I__4406 (
            .O(N__29521),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ));
    Odrv4 I__4405 (
            .O(N__29518),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ));
    InMux I__4404 (
            .O(N__29513),
            .I(N__29506));
    InMux I__4403 (
            .O(N__29512),
            .I(N__29506));
    InMux I__4402 (
            .O(N__29511),
            .I(N__29503));
    LocalMux I__4401 (
            .O(N__29506),
            .I(N__29500));
    LocalMux I__4400 (
            .O(N__29503),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ));
    Odrv4 I__4399 (
            .O(N__29500),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ));
    CascadeMux I__4398 (
            .O(N__29495),
            .I(N__29492));
    InMux I__4397 (
            .O(N__29492),
            .I(N__29487));
    InMux I__4396 (
            .O(N__29491),
            .I(N__29484));
    InMux I__4395 (
            .O(N__29490),
            .I(N__29481));
    LocalMux I__4394 (
            .O(N__29487),
            .I(N__29476));
    LocalMux I__4393 (
            .O(N__29484),
            .I(N__29476));
    LocalMux I__4392 (
            .O(N__29481),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ));
    Odrv12 I__4391 (
            .O(N__29476),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ));
    CascadeMux I__4390 (
            .O(N__29471),
            .I(N__29468));
    InMux I__4389 (
            .O(N__29468),
            .I(N__29464));
    InMux I__4388 (
            .O(N__29467),
            .I(N__29460));
    LocalMux I__4387 (
            .O(N__29464),
            .I(N__29457));
    InMux I__4386 (
            .O(N__29463),
            .I(N__29454));
    LocalMux I__4385 (
            .O(N__29460),
            .I(N__29451));
    Span4Mux_v I__4384 (
            .O(N__29457),
            .I(N__29448));
    LocalMux I__4383 (
            .O(N__29454),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ));
    Odrv4 I__4382 (
            .O(N__29451),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ));
    Odrv4 I__4381 (
            .O(N__29448),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ));
    InMux I__4380 (
            .O(N__29441),
            .I(N__29434));
    InMux I__4379 (
            .O(N__29440),
            .I(N__29434));
    InMux I__4378 (
            .O(N__29439),
            .I(N__29431));
    LocalMux I__4377 (
            .O(N__29434),
            .I(N__29428));
    LocalMux I__4376 (
            .O(N__29431),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ));
    Odrv12 I__4375 (
            .O(N__29428),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ));
    CascadeMux I__4374 (
            .O(N__29423),
            .I(N__29419));
    CascadeMux I__4373 (
            .O(N__29422),
            .I(N__29416));
    InMux I__4372 (
            .O(N__29419),
            .I(N__29410));
    InMux I__4371 (
            .O(N__29416),
            .I(N__29410));
    InMux I__4370 (
            .O(N__29415),
            .I(N__29407));
    LocalMux I__4369 (
            .O(N__29410),
            .I(N__29404));
    LocalMux I__4368 (
            .O(N__29407),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ));
    Odrv12 I__4367 (
            .O(N__29404),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ));
    InMux I__4366 (
            .O(N__29399),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_28 ));
    InMux I__4365 (
            .O(N__29396),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_29 ));
    InMux I__4364 (
            .O(N__29393),
            .I(N__29369));
    InMux I__4363 (
            .O(N__29392),
            .I(N__29369));
    InMux I__4362 (
            .O(N__29391),
            .I(N__29369));
    InMux I__4361 (
            .O(N__29390),
            .I(N__29369));
    InMux I__4360 (
            .O(N__29389),
            .I(N__29360));
    InMux I__4359 (
            .O(N__29388),
            .I(N__29360));
    InMux I__4358 (
            .O(N__29387),
            .I(N__29360));
    InMux I__4357 (
            .O(N__29386),
            .I(N__29360));
    InMux I__4356 (
            .O(N__29385),
            .I(N__29337));
    InMux I__4355 (
            .O(N__29384),
            .I(N__29337));
    InMux I__4354 (
            .O(N__29383),
            .I(N__29337));
    InMux I__4353 (
            .O(N__29382),
            .I(N__29326));
    InMux I__4352 (
            .O(N__29381),
            .I(N__29326));
    InMux I__4351 (
            .O(N__29380),
            .I(N__29326));
    InMux I__4350 (
            .O(N__29379),
            .I(N__29326));
    InMux I__4349 (
            .O(N__29378),
            .I(N__29326));
    LocalMux I__4348 (
            .O(N__29369),
            .I(N__29323));
    LocalMux I__4347 (
            .O(N__29360),
            .I(N__29320));
    InMux I__4346 (
            .O(N__29359),
            .I(N__29311));
    InMux I__4345 (
            .O(N__29358),
            .I(N__29311));
    InMux I__4344 (
            .O(N__29357),
            .I(N__29311));
    InMux I__4343 (
            .O(N__29356),
            .I(N__29311));
    InMux I__4342 (
            .O(N__29355),
            .I(N__29302));
    InMux I__4341 (
            .O(N__29354),
            .I(N__29302));
    InMux I__4340 (
            .O(N__29353),
            .I(N__29302));
    InMux I__4339 (
            .O(N__29352),
            .I(N__29302));
    InMux I__4338 (
            .O(N__29351),
            .I(N__29293));
    InMux I__4337 (
            .O(N__29350),
            .I(N__29293));
    InMux I__4336 (
            .O(N__29349),
            .I(N__29293));
    InMux I__4335 (
            .O(N__29348),
            .I(N__29293));
    InMux I__4334 (
            .O(N__29347),
            .I(N__29284));
    InMux I__4333 (
            .O(N__29346),
            .I(N__29284));
    InMux I__4332 (
            .O(N__29345),
            .I(N__29284));
    InMux I__4331 (
            .O(N__29344),
            .I(N__29284));
    LocalMux I__4330 (
            .O(N__29337),
            .I(N__29279));
    LocalMux I__4329 (
            .O(N__29326),
            .I(N__29279));
    Odrv4 I__4328 (
            .O(N__29323),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    Odrv4 I__4327 (
            .O(N__29320),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    LocalMux I__4326 (
            .O(N__29311),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    LocalMux I__4325 (
            .O(N__29302),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    LocalMux I__4324 (
            .O(N__29293),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    LocalMux I__4323 (
            .O(N__29284),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    Odrv4 I__4322 (
            .O(N__29279),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    InMux I__4321 (
            .O(N__29264),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_30 ));
    CEMux I__4320 (
            .O(N__29261),
            .I(N__29257));
    CEMux I__4319 (
            .O(N__29260),
            .I(N__29253));
    LocalMux I__4318 (
            .O(N__29257),
            .I(N__29250));
    CEMux I__4317 (
            .O(N__29256),
            .I(N__29246));
    LocalMux I__4316 (
            .O(N__29253),
            .I(N__29241));
    Span4Mux_v I__4315 (
            .O(N__29250),
            .I(N__29241));
    CEMux I__4314 (
            .O(N__29249),
            .I(N__29238));
    LocalMux I__4313 (
            .O(N__29246),
            .I(N__29233));
    Span4Mux_s1_v I__4312 (
            .O(N__29241),
            .I(N__29233));
    LocalMux I__4311 (
            .O(N__29238),
            .I(N__29230));
    Odrv4 I__4310 (
            .O(N__29233),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__4309 (
            .O(N__29230),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__4308 (
            .O(N__29225),
            .I(N__29220));
    InMux I__4307 (
            .O(N__29224),
            .I(N__29215));
    InMux I__4306 (
            .O(N__29223),
            .I(N__29215));
    LocalMux I__4305 (
            .O(N__29220),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ));
    LocalMux I__4304 (
            .O(N__29215),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ));
    InMux I__4303 (
            .O(N__29210),
            .I(N__29205));
    InMux I__4302 (
            .O(N__29209),
            .I(N__29200));
    InMux I__4301 (
            .O(N__29208),
            .I(N__29200));
    LocalMux I__4300 (
            .O(N__29205),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ));
    LocalMux I__4299 (
            .O(N__29200),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ));
    InMux I__4298 (
            .O(N__29195),
            .I(N__29190));
    InMux I__4297 (
            .O(N__29194),
            .I(N__29185));
    InMux I__4296 (
            .O(N__29193),
            .I(N__29185));
    LocalMux I__4295 (
            .O(N__29190),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ));
    LocalMux I__4294 (
            .O(N__29185),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ));
    InMux I__4293 (
            .O(N__29180),
            .I(N__29175));
    InMux I__4292 (
            .O(N__29179),
            .I(N__29172));
    InMux I__4291 (
            .O(N__29178),
            .I(N__29169));
    LocalMux I__4290 (
            .O(N__29175),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ));
    LocalMux I__4289 (
            .O(N__29172),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ));
    LocalMux I__4288 (
            .O(N__29169),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ));
    InMux I__4287 (
            .O(N__29162),
            .I(N__29155));
    InMux I__4286 (
            .O(N__29161),
            .I(N__29155));
    InMux I__4285 (
            .O(N__29160),
            .I(N__29152));
    LocalMux I__4284 (
            .O(N__29155),
            .I(N__29149));
    LocalMux I__4283 (
            .O(N__29152),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ));
    Odrv4 I__4282 (
            .O(N__29149),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ));
    CascadeMux I__4281 (
            .O(N__29144),
            .I(N__29140));
    CascadeMux I__4280 (
            .O(N__29143),
            .I(N__29137));
    InMux I__4279 (
            .O(N__29140),
            .I(N__29131));
    InMux I__4278 (
            .O(N__29137),
            .I(N__29131));
    InMux I__4277 (
            .O(N__29136),
            .I(N__29128));
    LocalMux I__4276 (
            .O(N__29131),
            .I(N__29125));
    LocalMux I__4275 (
            .O(N__29128),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ));
    Odrv4 I__4274 (
            .O(N__29125),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ));
    InMux I__4273 (
            .O(N__29120),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_19 ));
    InMux I__4272 (
            .O(N__29117),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_20 ));
    InMux I__4271 (
            .O(N__29114),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_21 ));
    InMux I__4270 (
            .O(N__29111),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_22 ));
    InMux I__4269 (
            .O(N__29108),
            .I(bfn_10_5_0_));
    InMux I__4268 (
            .O(N__29105),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_24 ));
    InMux I__4267 (
            .O(N__29102),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_25 ));
    InMux I__4266 (
            .O(N__29099),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_26 ));
    InMux I__4265 (
            .O(N__29096),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_27 ));
    InMux I__4264 (
            .O(N__29093),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_10 ));
    InMux I__4263 (
            .O(N__29090),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_11 ));
    InMux I__4262 (
            .O(N__29087),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_12 ));
    InMux I__4261 (
            .O(N__29084),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_13 ));
    InMux I__4260 (
            .O(N__29081),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_14 ));
    InMux I__4259 (
            .O(N__29078),
            .I(bfn_10_4_0_));
    InMux I__4258 (
            .O(N__29075),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_16 ));
    InMux I__4257 (
            .O(N__29072),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_17 ));
    InMux I__4256 (
            .O(N__29069),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_18 ));
    InMux I__4255 (
            .O(N__29066),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_1 ));
    InMux I__4254 (
            .O(N__29063),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_2 ));
    InMux I__4253 (
            .O(N__29060),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_3 ));
    InMux I__4252 (
            .O(N__29057),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_4 ));
    InMux I__4251 (
            .O(N__29054),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_5 ));
    InMux I__4250 (
            .O(N__29051),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_6 ));
    InMux I__4249 (
            .O(N__29048),
            .I(bfn_10_3_0_));
    InMux I__4248 (
            .O(N__29045),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_8 ));
    InMux I__4247 (
            .O(N__29042),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_9 ));
    InMux I__4246 (
            .O(N__29039),
            .I(N__29036));
    LocalMux I__4245 (
            .O(N__29036),
            .I(N__29033));
    Odrv4 I__4244 (
            .O(N__29033),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ));
    InMux I__4243 (
            .O(N__29030),
            .I(N__29027));
    LocalMux I__4242 (
            .O(N__29027),
            .I(N__29023));
    CascadeMux I__4241 (
            .O(N__29026),
            .I(N__29020));
    Span12Mux_s10_h I__4240 (
            .O(N__29023),
            .I(N__29016));
    InMux I__4239 (
            .O(N__29020),
            .I(N__29011));
    InMux I__4238 (
            .O(N__29019),
            .I(N__29011));
    Span12Mux_v I__4237 (
            .O(N__29016),
            .I(N__29008));
    LocalMux I__4236 (
            .O(N__29011),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    Odrv12 I__4235 (
            .O(N__29008),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    IoInMux I__4234 (
            .O(N__29003),
            .I(N__29000));
    LocalMux I__4233 (
            .O(N__29000),
            .I(N__28997));
    Span4Mux_s3_v I__4232 (
            .O(N__28997),
            .I(N__28994));
    Span4Mux_v I__4231 (
            .O(N__28994),
            .I(N__28991));
    Odrv4 I__4230 (
            .O(N__28991),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__4229 (
            .O(N__28988),
            .I(N__28983));
    InMux I__4228 (
            .O(N__28987),
            .I(N__28978));
    InMux I__4227 (
            .O(N__28986),
            .I(N__28978));
    LocalMux I__4226 (
            .O(N__28983),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ));
    LocalMux I__4225 (
            .O(N__28978),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ));
    CascadeMux I__4224 (
            .O(N__28973),
            .I(N__28969));
    InMux I__4223 (
            .O(N__28972),
            .I(N__28962));
    InMux I__4222 (
            .O(N__28969),
            .I(N__28962));
    InMux I__4221 (
            .O(N__28968),
            .I(N__28957));
    InMux I__4220 (
            .O(N__28967),
            .I(N__28957));
    LocalMux I__4219 (
            .O(N__28962),
            .I(N__28954));
    LocalMux I__4218 (
            .O(N__28957),
            .I(N__28949));
    Span12Mux_s8_v I__4217 (
            .O(N__28954),
            .I(N__28949));
    Span12Mux_v I__4216 (
            .O(N__28949),
            .I(N__28946));
    Odrv12 I__4215 (
            .O(N__28946),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ));
    InMux I__4214 (
            .O(N__28943),
            .I(N__28938));
    InMux I__4213 (
            .O(N__28942),
            .I(N__28933));
    InMux I__4212 (
            .O(N__28941),
            .I(N__28933));
    LocalMux I__4211 (
            .O(N__28938),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ));
    LocalMux I__4210 (
            .O(N__28933),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ));
    CascadeMux I__4209 (
            .O(N__28928),
            .I(N__28925));
    InMux I__4208 (
            .O(N__28925),
            .I(N__28922));
    LocalMux I__4207 (
            .O(N__28922),
            .I(N__28919));
    Odrv4 I__4206 (
            .O(N__28919),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt30 ));
    CascadeMux I__4205 (
            .O(N__28916),
            .I(N__28913));
    InMux I__4204 (
            .O(N__28913),
            .I(N__28909));
    InMux I__4203 (
            .O(N__28912),
            .I(N__28905));
    LocalMux I__4202 (
            .O(N__28909),
            .I(N__28902));
    InMux I__4201 (
            .O(N__28908),
            .I(N__28899));
    LocalMux I__4200 (
            .O(N__28905),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ));
    Odrv4 I__4199 (
            .O(N__28902),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ));
    LocalMux I__4198 (
            .O(N__28899),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ));
    InMux I__4197 (
            .O(N__28892),
            .I(N__28888));
    InMux I__4196 (
            .O(N__28891),
            .I(N__28885));
    LocalMux I__4195 (
            .O(N__28888),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ));
    LocalMux I__4194 (
            .O(N__28885),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ));
    CascadeMux I__4193 (
            .O(N__28880),
            .I(N__28875));
    InMux I__4192 (
            .O(N__28879),
            .I(N__28872));
    InMux I__4191 (
            .O(N__28878),
            .I(N__28867));
    InMux I__4190 (
            .O(N__28875),
            .I(N__28867));
    LocalMux I__4189 (
            .O(N__28872),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ));
    LocalMux I__4188 (
            .O(N__28867),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ));
    InMux I__4187 (
            .O(N__28862),
            .I(N__28856));
    InMux I__4186 (
            .O(N__28861),
            .I(N__28856));
    LocalMux I__4185 (
            .O(N__28856),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ));
    CascadeMux I__4184 (
            .O(N__28853),
            .I(N__28850));
    InMux I__4183 (
            .O(N__28850),
            .I(N__28847));
    LocalMux I__4182 (
            .O(N__28847),
            .I(N__28844));
    Span4Mux_h I__4181 (
            .O(N__28844),
            .I(N__28841));
    Odrv4 I__4180 (
            .O(N__28841),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt24 ));
    InMux I__4179 (
            .O(N__28838),
            .I(N__28818));
    InMux I__4178 (
            .O(N__28837),
            .I(N__28818));
    InMux I__4177 (
            .O(N__28836),
            .I(N__28818));
    InMux I__4176 (
            .O(N__28835),
            .I(N__28818));
    InMux I__4175 (
            .O(N__28834),
            .I(N__28797));
    InMux I__4174 (
            .O(N__28833),
            .I(N__28797));
    InMux I__4173 (
            .O(N__28832),
            .I(N__28797));
    InMux I__4172 (
            .O(N__28831),
            .I(N__28797));
    InMux I__4171 (
            .O(N__28830),
            .I(N__28788));
    InMux I__4170 (
            .O(N__28829),
            .I(N__28788));
    InMux I__4169 (
            .O(N__28828),
            .I(N__28788));
    InMux I__4168 (
            .O(N__28827),
            .I(N__28788));
    LocalMux I__4167 (
            .O(N__28818),
            .I(N__28777));
    InMux I__4166 (
            .O(N__28817),
            .I(N__28768));
    InMux I__4165 (
            .O(N__28816),
            .I(N__28768));
    InMux I__4164 (
            .O(N__28815),
            .I(N__28768));
    InMux I__4163 (
            .O(N__28814),
            .I(N__28768));
    InMux I__4162 (
            .O(N__28813),
            .I(N__28759));
    InMux I__4161 (
            .O(N__28812),
            .I(N__28759));
    InMux I__4160 (
            .O(N__28811),
            .I(N__28759));
    InMux I__4159 (
            .O(N__28810),
            .I(N__28759));
    InMux I__4158 (
            .O(N__28809),
            .I(N__28750));
    InMux I__4157 (
            .O(N__28808),
            .I(N__28750));
    InMux I__4156 (
            .O(N__28807),
            .I(N__28750));
    InMux I__4155 (
            .O(N__28806),
            .I(N__28750));
    LocalMux I__4154 (
            .O(N__28797),
            .I(N__28745));
    LocalMux I__4153 (
            .O(N__28788),
            .I(N__28745));
    InMux I__4152 (
            .O(N__28787),
            .I(N__28736));
    InMux I__4151 (
            .O(N__28786),
            .I(N__28736));
    InMux I__4150 (
            .O(N__28785),
            .I(N__28736));
    InMux I__4149 (
            .O(N__28784),
            .I(N__28736));
    InMux I__4148 (
            .O(N__28783),
            .I(N__28727));
    InMux I__4147 (
            .O(N__28782),
            .I(N__28727));
    InMux I__4146 (
            .O(N__28781),
            .I(N__28727));
    InMux I__4145 (
            .O(N__28780),
            .I(N__28727));
    Span4Mux_h I__4144 (
            .O(N__28777),
            .I(N__28722));
    LocalMux I__4143 (
            .O(N__28768),
            .I(N__28722));
    LocalMux I__4142 (
            .O(N__28759),
            .I(N__28715));
    LocalMux I__4141 (
            .O(N__28750),
            .I(N__28715));
    Span4Mux_h I__4140 (
            .O(N__28745),
            .I(N__28715));
    LocalMux I__4139 (
            .O(N__28736),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    LocalMux I__4138 (
            .O(N__28727),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    Odrv4 I__4137 (
            .O(N__28722),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    Odrv4 I__4136 (
            .O(N__28715),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    InMux I__4135 (
            .O(N__28706),
            .I(N__28703));
    LocalMux I__4134 (
            .O(N__28703),
            .I(N__28700));
    Span4Mux_h I__4133 (
            .O(N__28700),
            .I(N__28696));
    CascadeMux I__4132 (
            .O(N__28699),
            .I(N__28692));
    Sp12to4 I__4131 (
            .O(N__28696),
            .I(N__28688));
    InMux I__4130 (
            .O(N__28695),
            .I(N__28683));
    InMux I__4129 (
            .O(N__28692),
            .I(N__28683));
    InMux I__4128 (
            .O(N__28691),
            .I(N__28680));
    Span12Mux_v I__4127 (
            .O(N__28688),
            .I(N__28677));
    LocalMux I__4126 (
            .O(N__28683),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__4125 (
            .O(N__28680),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__4124 (
            .O(N__28677),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    IoInMux I__4123 (
            .O(N__28670),
            .I(N__28667));
    LocalMux I__4122 (
            .O(N__28667),
            .I(N__28664));
    Odrv4 I__4121 (
            .O(N__28664),
            .I(s3_phy_c));
    InMux I__4120 (
            .O(N__28661),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_0 ));
    InMux I__4119 (
            .O(N__28658),
            .I(N__28655));
    LocalMux I__4118 (
            .O(N__28655),
            .I(N__28652));
    Span4Mux_h I__4117 (
            .O(N__28652),
            .I(N__28648));
    InMux I__4116 (
            .O(N__28651),
            .I(N__28645));
    Odrv4 I__4115 (
            .O(N__28648),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ));
    LocalMux I__4114 (
            .O(N__28645),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ));
    InMux I__4113 (
            .O(N__28640),
            .I(N__28635));
    InMux I__4112 (
            .O(N__28639),
            .I(N__28632));
    InMux I__4111 (
            .O(N__28638),
            .I(N__28629));
    LocalMux I__4110 (
            .O(N__28635),
            .I(N__28626));
    LocalMux I__4109 (
            .O(N__28632),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ));
    LocalMux I__4108 (
            .O(N__28629),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ));
    Odrv4 I__4107 (
            .O(N__28626),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ));
    CascadeMux I__4106 (
            .O(N__28619),
            .I(N__28615));
    CascadeMux I__4105 (
            .O(N__28618),
            .I(N__28611));
    InMux I__4104 (
            .O(N__28615),
            .I(N__28608));
    InMux I__4103 (
            .O(N__28614),
            .I(N__28605));
    InMux I__4102 (
            .O(N__28611),
            .I(N__28602));
    LocalMux I__4101 (
            .O(N__28608),
            .I(N__28599));
    LocalMux I__4100 (
            .O(N__28605),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ));
    LocalMux I__4099 (
            .O(N__28602),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ));
    Odrv4 I__4098 (
            .O(N__28599),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ));
    InMux I__4097 (
            .O(N__28592),
            .I(N__28589));
    LocalMux I__4096 (
            .O(N__28589),
            .I(N__28586));
    Span4Mux_h I__4095 (
            .O(N__28586),
            .I(N__28582));
    InMux I__4094 (
            .O(N__28585),
            .I(N__28579));
    Odrv4 I__4093 (
            .O(N__28582),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ));
    LocalMux I__4092 (
            .O(N__28579),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ));
    InMux I__4091 (
            .O(N__28574),
            .I(N__28571));
    LocalMux I__4090 (
            .O(N__28571),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt16 ));
    InMux I__4089 (
            .O(N__28568),
            .I(N__28562));
    InMux I__4088 (
            .O(N__28567),
            .I(N__28562));
    LocalMux I__4087 (
            .O(N__28562),
            .I(N__28558));
    InMux I__4086 (
            .O(N__28561),
            .I(N__28555));
    Span4Mux_h I__4085 (
            .O(N__28558),
            .I(N__28552));
    LocalMux I__4084 (
            .O(N__28555),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ));
    Odrv4 I__4083 (
            .O(N__28552),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ));
    InMux I__4082 (
            .O(N__28547),
            .I(N__28540));
    InMux I__4081 (
            .O(N__28546),
            .I(N__28540));
    InMux I__4080 (
            .O(N__28545),
            .I(N__28537));
    LocalMux I__4079 (
            .O(N__28540),
            .I(N__28534));
    LocalMux I__4078 (
            .O(N__28537),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ));
    Odrv4 I__4077 (
            .O(N__28534),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ));
    InMux I__4076 (
            .O(N__28529),
            .I(N__28526));
    LocalMux I__4075 (
            .O(N__28526),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt28 ));
    InMux I__4074 (
            .O(N__28523),
            .I(N__28520));
    LocalMux I__4073 (
            .O(N__28520),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ));
    InMux I__4072 (
            .O(N__28517),
            .I(N__28514));
    LocalMux I__4071 (
            .O(N__28514),
            .I(N__28511));
    Span4Mux_v I__4070 (
            .O(N__28511),
            .I(N__28507));
    InMux I__4069 (
            .O(N__28510),
            .I(N__28504));
    Odrv4 I__4068 (
            .O(N__28507),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_24));
    LocalMux I__4067 (
            .O(N__28504),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_24));
    InMux I__4066 (
            .O(N__28499),
            .I(N__28495));
    InMux I__4065 (
            .O(N__28498),
            .I(N__28492));
    LocalMux I__4064 (
            .O(N__28495),
            .I(N__28489));
    LocalMux I__4063 (
            .O(N__28492),
            .I(N__28486));
    Span4Mux_v I__4062 (
            .O(N__28489),
            .I(N__28481));
    Span4Mux_v I__4061 (
            .O(N__28486),
            .I(N__28481));
    Odrv4 I__4060 (
            .O(N__28481),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_25));
    InMux I__4059 (
            .O(N__28478),
            .I(N__28475));
    LocalMux I__4058 (
            .O(N__28475),
            .I(N__28472));
    Odrv4 I__4057 (
            .O(N__28472),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt26 ));
    InMux I__4056 (
            .O(N__28469),
            .I(N__28466));
    LocalMux I__4055 (
            .O(N__28466),
            .I(N__28462));
    InMux I__4054 (
            .O(N__28465),
            .I(N__28459));
    Span4Mux_h I__4053 (
            .O(N__28462),
            .I(N__28456));
    LocalMux I__4052 (
            .O(N__28459),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_26));
    Odrv4 I__4051 (
            .O(N__28456),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_26));
    InMux I__4050 (
            .O(N__28451),
            .I(N__28446));
    InMux I__4049 (
            .O(N__28450),
            .I(N__28441));
    InMux I__4048 (
            .O(N__28449),
            .I(N__28441));
    LocalMux I__4047 (
            .O(N__28446),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ));
    LocalMux I__4046 (
            .O(N__28441),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ));
    InMux I__4045 (
            .O(N__28436),
            .I(N__28430));
    InMux I__4044 (
            .O(N__28435),
            .I(N__28430));
    LocalMux I__4043 (
            .O(N__28430),
            .I(N__28427));
    Odrv4 I__4042 (
            .O(N__28427),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ));
    CascadeMux I__4041 (
            .O(N__28424),
            .I(N__28420));
    CascadeMux I__4040 (
            .O(N__28423),
            .I(N__28417));
    InMux I__4039 (
            .O(N__28420),
            .I(N__28412));
    InMux I__4038 (
            .O(N__28417),
            .I(N__28412));
    LocalMux I__4037 (
            .O(N__28412),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ));
    InMux I__4036 (
            .O(N__28409),
            .I(N__28404));
    InMux I__4035 (
            .O(N__28408),
            .I(N__28399));
    InMux I__4034 (
            .O(N__28407),
            .I(N__28399));
    LocalMux I__4033 (
            .O(N__28404),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ));
    LocalMux I__4032 (
            .O(N__28399),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ));
    CascadeMux I__4031 (
            .O(N__28394),
            .I(N__28391));
    InMux I__4030 (
            .O(N__28391),
            .I(N__28388));
    LocalMux I__4029 (
            .O(N__28388),
            .I(N__28385));
    Odrv4 I__4028 (
            .O(N__28385),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ));
    InMux I__4027 (
            .O(N__28382),
            .I(N__28379));
    LocalMux I__4026 (
            .O(N__28379),
            .I(N__28376));
    Odrv4 I__4025 (
            .O(N__28376),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ));
    InMux I__4024 (
            .O(N__28373),
            .I(bfn_9_21_0_));
    InMux I__4023 (
            .O(N__28370),
            .I(N__28364));
    InMux I__4022 (
            .O(N__28369),
            .I(N__28364));
    LocalMux I__4021 (
            .O(N__28364),
            .I(N__28360));
    InMux I__4020 (
            .O(N__28363),
            .I(N__28357));
    Odrv12 I__4019 (
            .O(N__28360),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ));
    LocalMux I__4018 (
            .O(N__28357),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ));
    CascadeMux I__4017 (
            .O(N__28352),
            .I(N__28348));
    InMux I__4016 (
            .O(N__28351),
            .I(N__28345));
    InMux I__4015 (
            .O(N__28348),
            .I(N__28342));
    LocalMux I__4014 (
            .O(N__28345),
            .I(\phase_controller_inst1.stoper_tr.counter ));
    LocalMux I__4013 (
            .O(N__28342),
            .I(\phase_controller_inst1.stoper_tr.counter ));
    CascadeMux I__4012 (
            .O(N__28337),
            .I(N__28334));
    InMux I__4011 (
            .O(N__28334),
            .I(N__28331));
    LocalMux I__4010 (
            .O(N__28331),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ));
    InMux I__4009 (
            .O(N__28328),
            .I(N__28325));
    LocalMux I__4008 (
            .O(N__28325),
            .I(N__28322));
    Span4Mux_v I__4007 (
            .O(N__28322),
            .I(N__28319));
    Odrv4 I__4006 (
            .O(N__28319),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ));
    InMux I__4005 (
            .O(N__28316),
            .I(N__28312));
    InMux I__4004 (
            .O(N__28315),
            .I(N__28309));
    LocalMux I__4003 (
            .O(N__28312),
            .I(N__28306));
    LocalMux I__4002 (
            .O(N__28309),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ));
    Odrv4 I__4001 (
            .O(N__28306),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ));
    CascadeMux I__4000 (
            .O(N__28301),
            .I(N__28298));
    InMux I__3999 (
            .O(N__28298),
            .I(N__28295));
    LocalMux I__3998 (
            .O(N__28295),
            .I(\phase_controller_inst1.stoper_tr.counter_i_11 ));
    CascadeMux I__3997 (
            .O(N__28292),
            .I(N__28289));
    InMux I__3996 (
            .O(N__28289),
            .I(N__28286));
    LocalMux I__3995 (
            .O(N__28286),
            .I(N__28283));
    Span4Mux_v I__3994 (
            .O(N__28283),
            .I(N__28280));
    Odrv4 I__3993 (
            .O(N__28280),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ));
    InMux I__3992 (
            .O(N__28277),
            .I(N__28273));
    InMux I__3991 (
            .O(N__28276),
            .I(N__28270));
    LocalMux I__3990 (
            .O(N__28273),
            .I(N__28267));
    LocalMux I__3989 (
            .O(N__28270),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ));
    Odrv4 I__3988 (
            .O(N__28267),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ));
    InMux I__3987 (
            .O(N__28262),
            .I(N__28259));
    LocalMux I__3986 (
            .O(N__28259),
            .I(\phase_controller_inst1.stoper_tr.counter_i_12 ));
    InMux I__3985 (
            .O(N__28256),
            .I(N__28252));
    InMux I__3984 (
            .O(N__28255),
            .I(N__28249));
    LocalMux I__3983 (
            .O(N__28252),
            .I(N__28246));
    LocalMux I__3982 (
            .O(N__28249),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ));
    Odrv4 I__3981 (
            .O(N__28246),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ));
    InMux I__3980 (
            .O(N__28241),
            .I(N__28238));
    LocalMux I__3979 (
            .O(N__28238),
            .I(N__28235));
    Span4Mux_v I__3978 (
            .O(N__28235),
            .I(N__28232));
    Odrv4 I__3977 (
            .O(N__28232),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ));
    CascadeMux I__3976 (
            .O(N__28229),
            .I(N__28226));
    InMux I__3975 (
            .O(N__28226),
            .I(N__28223));
    LocalMux I__3974 (
            .O(N__28223),
            .I(\phase_controller_inst1.stoper_tr.counter_i_13 ));
    InMux I__3973 (
            .O(N__28220),
            .I(N__28216));
    InMux I__3972 (
            .O(N__28219),
            .I(N__28213));
    LocalMux I__3971 (
            .O(N__28216),
            .I(N__28210));
    LocalMux I__3970 (
            .O(N__28213),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ));
    Odrv4 I__3969 (
            .O(N__28210),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ));
    InMux I__3968 (
            .O(N__28205),
            .I(N__28202));
    LocalMux I__3967 (
            .O(N__28202),
            .I(N__28199));
    Span4Mux_h I__3966 (
            .O(N__28199),
            .I(N__28196));
    Odrv4 I__3965 (
            .O(N__28196),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ));
    CascadeMux I__3964 (
            .O(N__28193),
            .I(N__28190));
    InMux I__3963 (
            .O(N__28190),
            .I(N__28187));
    LocalMux I__3962 (
            .O(N__28187),
            .I(\phase_controller_inst1.stoper_tr.counter_i_14 ));
    InMux I__3961 (
            .O(N__28184),
            .I(N__28180));
    InMux I__3960 (
            .O(N__28183),
            .I(N__28177));
    LocalMux I__3959 (
            .O(N__28180),
            .I(N__28174));
    LocalMux I__3958 (
            .O(N__28177),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ));
    Odrv4 I__3957 (
            .O(N__28174),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ));
    InMux I__3956 (
            .O(N__28169),
            .I(N__28166));
    LocalMux I__3955 (
            .O(N__28166),
            .I(N__28163));
    Span4Mux_h I__3954 (
            .O(N__28163),
            .I(N__28160));
    Odrv4 I__3953 (
            .O(N__28160),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ));
    CascadeMux I__3952 (
            .O(N__28157),
            .I(N__28154));
    InMux I__3951 (
            .O(N__28154),
            .I(N__28151));
    LocalMux I__3950 (
            .O(N__28151),
            .I(\phase_controller_inst1.stoper_tr.counter_i_15 ));
    CascadeMux I__3949 (
            .O(N__28148),
            .I(N__28145));
    InMux I__3948 (
            .O(N__28145),
            .I(N__28142));
    LocalMux I__3947 (
            .O(N__28142),
            .I(N__28139));
    Span4Mux_h I__3946 (
            .O(N__28139),
            .I(N__28136));
    Odrv4 I__3945 (
            .O(N__28136),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ));
    InMux I__3944 (
            .O(N__28133),
            .I(N__28130));
    LocalMux I__3943 (
            .O(N__28130),
            .I(N__28127));
    Odrv12 I__3942 (
            .O(N__28127),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ));
    CascadeMux I__3941 (
            .O(N__28124),
            .I(N__28121));
    InMux I__3940 (
            .O(N__28121),
            .I(N__28118));
    LocalMux I__3939 (
            .O(N__28118),
            .I(N__28115));
    Odrv4 I__3938 (
            .O(N__28115),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt18 ));
    CascadeMux I__3937 (
            .O(N__28112),
            .I(N__28109));
    InMux I__3936 (
            .O(N__28109),
            .I(N__28106));
    LocalMux I__3935 (
            .O(N__28106),
            .I(\phase_controller_inst1.stoper_tr.counter_i_3 ));
    InMux I__3934 (
            .O(N__28103),
            .I(N__28100));
    LocalMux I__3933 (
            .O(N__28100),
            .I(N__28097));
    Odrv12 I__3932 (
            .O(N__28097),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ));
    InMux I__3931 (
            .O(N__28094),
            .I(N__28090));
    InMux I__3930 (
            .O(N__28093),
            .I(N__28087));
    LocalMux I__3929 (
            .O(N__28090),
            .I(N__28084));
    LocalMux I__3928 (
            .O(N__28087),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ));
    Odrv4 I__3927 (
            .O(N__28084),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ));
    CascadeMux I__3926 (
            .O(N__28079),
            .I(N__28076));
    InMux I__3925 (
            .O(N__28076),
            .I(N__28073));
    LocalMux I__3924 (
            .O(N__28073),
            .I(N__28070));
    Odrv4 I__3923 (
            .O(N__28070),
            .I(\phase_controller_inst1.stoper_tr.counter_i_4 ));
    InMux I__3922 (
            .O(N__28067),
            .I(N__28063));
    InMux I__3921 (
            .O(N__28066),
            .I(N__28060));
    LocalMux I__3920 (
            .O(N__28063),
            .I(N__28057));
    LocalMux I__3919 (
            .O(N__28060),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ));
    Odrv4 I__3918 (
            .O(N__28057),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ));
    InMux I__3917 (
            .O(N__28052),
            .I(N__28049));
    LocalMux I__3916 (
            .O(N__28049),
            .I(N__28046));
    Odrv4 I__3915 (
            .O(N__28046),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ));
    CascadeMux I__3914 (
            .O(N__28043),
            .I(N__28040));
    InMux I__3913 (
            .O(N__28040),
            .I(N__28037));
    LocalMux I__3912 (
            .O(N__28037),
            .I(\phase_controller_inst1.stoper_tr.counter_i_5 ));
    InMux I__3911 (
            .O(N__28034),
            .I(N__28030));
    InMux I__3910 (
            .O(N__28033),
            .I(N__28027));
    LocalMux I__3909 (
            .O(N__28030),
            .I(N__28024));
    LocalMux I__3908 (
            .O(N__28027),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ));
    Odrv4 I__3907 (
            .O(N__28024),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ));
    InMux I__3906 (
            .O(N__28019),
            .I(N__28016));
    LocalMux I__3905 (
            .O(N__28016),
            .I(N__28013));
    Odrv12 I__3904 (
            .O(N__28013),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ));
    CascadeMux I__3903 (
            .O(N__28010),
            .I(N__28007));
    InMux I__3902 (
            .O(N__28007),
            .I(N__28004));
    LocalMux I__3901 (
            .O(N__28004),
            .I(\phase_controller_inst1.stoper_tr.counter_i_6 ));
    InMux I__3900 (
            .O(N__28001),
            .I(N__27998));
    LocalMux I__3899 (
            .O(N__27998),
            .I(N__27994));
    InMux I__3898 (
            .O(N__27997),
            .I(N__27991));
    Span4Mux_v I__3897 (
            .O(N__27994),
            .I(N__27988));
    LocalMux I__3896 (
            .O(N__27991),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ));
    Odrv4 I__3895 (
            .O(N__27988),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ));
    InMux I__3894 (
            .O(N__27983),
            .I(N__27980));
    LocalMux I__3893 (
            .O(N__27980),
            .I(N__27977));
    Odrv4 I__3892 (
            .O(N__27977),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ));
    CascadeMux I__3891 (
            .O(N__27974),
            .I(N__27971));
    InMux I__3890 (
            .O(N__27971),
            .I(N__27968));
    LocalMux I__3889 (
            .O(N__27968),
            .I(\phase_controller_inst1.stoper_tr.counter_i_7 ));
    CascadeMux I__3888 (
            .O(N__27965),
            .I(N__27962));
    InMux I__3887 (
            .O(N__27962),
            .I(N__27959));
    LocalMux I__3886 (
            .O(N__27959),
            .I(N__27956));
    Span4Mux_v I__3885 (
            .O(N__27956),
            .I(N__27953));
    Odrv4 I__3884 (
            .O(N__27953),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ));
    InMux I__3883 (
            .O(N__27950),
            .I(N__27947));
    LocalMux I__3882 (
            .O(N__27947),
            .I(N__27943));
    InMux I__3881 (
            .O(N__27946),
            .I(N__27940));
    Span4Mux_h I__3880 (
            .O(N__27943),
            .I(N__27937));
    LocalMux I__3879 (
            .O(N__27940),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ));
    Odrv4 I__3878 (
            .O(N__27937),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ));
    InMux I__3877 (
            .O(N__27932),
            .I(N__27929));
    LocalMux I__3876 (
            .O(N__27929),
            .I(\phase_controller_inst1.stoper_tr.counter_i_8 ));
    InMux I__3875 (
            .O(N__27926),
            .I(N__27923));
    LocalMux I__3874 (
            .O(N__27923),
            .I(N__27920));
    Span4Mux_v I__3873 (
            .O(N__27920),
            .I(N__27917));
    Odrv4 I__3872 (
            .O(N__27917),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ));
    InMux I__3871 (
            .O(N__27914),
            .I(N__27910));
    InMux I__3870 (
            .O(N__27913),
            .I(N__27907));
    LocalMux I__3869 (
            .O(N__27910),
            .I(N__27904));
    LocalMux I__3868 (
            .O(N__27907),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ));
    Odrv4 I__3867 (
            .O(N__27904),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ));
    CascadeMux I__3866 (
            .O(N__27899),
            .I(N__27896));
    InMux I__3865 (
            .O(N__27896),
            .I(N__27893));
    LocalMux I__3864 (
            .O(N__27893),
            .I(\phase_controller_inst1.stoper_tr.counter_i_9 ));
    CascadeMux I__3863 (
            .O(N__27890),
            .I(N__27887));
    InMux I__3862 (
            .O(N__27887),
            .I(N__27884));
    LocalMux I__3861 (
            .O(N__27884),
            .I(N__27881));
    Span4Mux_v I__3860 (
            .O(N__27881),
            .I(N__27878));
    Odrv4 I__3859 (
            .O(N__27878),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ));
    InMux I__3858 (
            .O(N__27875),
            .I(N__27871));
    InMux I__3857 (
            .O(N__27874),
            .I(N__27868));
    LocalMux I__3856 (
            .O(N__27871),
            .I(N__27865));
    LocalMux I__3855 (
            .O(N__27868),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ));
    Odrv4 I__3854 (
            .O(N__27865),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ));
    InMux I__3853 (
            .O(N__27860),
            .I(N__27857));
    LocalMux I__3852 (
            .O(N__27857),
            .I(\phase_controller_inst1.stoper_tr.counter_i_10 ));
    InMux I__3851 (
            .O(N__27854),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ));
    InMux I__3850 (
            .O(N__27851),
            .I(N__27848));
    LocalMux I__3849 (
            .O(N__27848),
            .I(N__27844));
    InMux I__3848 (
            .O(N__27847),
            .I(N__27841));
    Span4Mux_h I__3847 (
            .O(N__27844),
            .I(N__27838));
    LocalMux I__3846 (
            .O(N__27841),
            .I(N__27835));
    Odrv4 I__3845 (
            .O(N__27838),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ));
    Odrv4 I__3844 (
            .O(N__27835),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ));
    InMux I__3843 (
            .O(N__27830),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ));
    InMux I__3842 (
            .O(N__27827),
            .I(N__27823));
    InMux I__3841 (
            .O(N__27826),
            .I(N__27820));
    LocalMux I__3840 (
            .O(N__27823),
            .I(N__27817));
    LocalMux I__3839 (
            .O(N__27820),
            .I(N__27812));
    Span4Mux_h I__3838 (
            .O(N__27817),
            .I(N__27812));
    Odrv4 I__3837 (
            .O(N__27812),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ));
    InMux I__3836 (
            .O(N__27809),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ));
    InMux I__3835 (
            .O(N__27806),
            .I(N__27803));
    LocalMux I__3834 (
            .O(N__27803),
            .I(N__27800));
    Odrv4 I__3833 (
            .O(N__27800),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ));
    InMux I__3832 (
            .O(N__27797),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ));
    InMux I__3831 (
            .O(N__27794),
            .I(N__27790));
    InMux I__3830 (
            .O(N__27793),
            .I(N__27787));
    LocalMux I__3829 (
            .O(N__27790),
            .I(N__27784));
    LocalMux I__3828 (
            .O(N__27787),
            .I(N__27781));
    Span4Mux_v I__3827 (
            .O(N__27784),
            .I(N__27778));
    Span4Mux_h I__3826 (
            .O(N__27781),
            .I(N__27775));
    Span4Mux_v I__3825 (
            .O(N__27778),
            .I(N__27772));
    Odrv4 I__3824 (
            .O(N__27775),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_28));
    Odrv4 I__3823 (
            .O(N__27772),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_28));
    InMux I__3822 (
            .O(N__27767),
            .I(N__27764));
    LocalMux I__3821 (
            .O(N__27764),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ));
    InMux I__3820 (
            .O(N__27761),
            .I(N__27758));
    LocalMux I__3819 (
            .O(N__27758),
            .I(N__27754));
    InMux I__3818 (
            .O(N__27757),
            .I(N__27751));
    Span4Mux_h I__3817 (
            .O(N__27754),
            .I(N__27748));
    LocalMux I__3816 (
            .O(N__27751),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ));
    Odrv4 I__3815 (
            .O(N__27748),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ));
    CascadeMux I__3814 (
            .O(N__27743),
            .I(N__27740));
    InMux I__3813 (
            .O(N__27740),
            .I(N__27737));
    LocalMux I__3812 (
            .O(N__27737),
            .I(\phase_controller_inst1.stoper_tr.counter_i_0 ));
    InMux I__3811 (
            .O(N__27734),
            .I(N__27731));
    LocalMux I__3810 (
            .O(N__27731),
            .I(N__27728));
    Span4Mux_v I__3809 (
            .O(N__27728),
            .I(N__27725));
    Odrv4 I__3808 (
            .O(N__27725),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ));
    InMux I__3807 (
            .O(N__27722),
            .I(N__27718));
    InMux I__3806 (
            .O(N__27721),
            .I(N__27715));
    LocalMux I__3805 (
            .O(N__27718),
            .I(N__27712));
    LocalMux I__3804 (
            .O(N__27715),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ));
    Odrv4 I__3803 (
            .O(N__27712),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ));
    CascadeMux I__3802 (
            .O(N__27707),
            .I(N__27704));
    InMux I__3801 (
            .O(N__27704),
            .I(N__27701));
    LocalMux I__3800 (
            .O(N__27701),
            .I(N__27698));
    Odrv4 I__3799 (
            .O(N__27698),
            .I(\phase_controller_inst1.stoper_tr.counter_i_1 ));
    InMux I__3798 (
            .O(N__27695),
            .I(N__27692));
    LocalMux I__3797 (
            .O(N__27692),
            .I(N__27689));
    Span4Mux_h I__3796 (
            .O(N__27689),
            .I(N__27686));
    Odrv4 I__3795 (
            .O(N__27686),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ));
    InMux I__3794 (
            .O(N__27683),
            .I(N__27679));
    InMux I__3793 (
            .O(N__27682),
            .I(N__27676));
    LocalMux I__3792 (
            .O(N__27679),
            .I(N__27673));
    LocalMux I__3791 (
            .O(N__27676),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ));
    Odrv4 I__3790 (
            .O(N__27673),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ));
    CascadeMux I__3789 (
            .O(N__27668),
            .I(N__27665));
    InMux I__3788 (
            .O(N__27665),
            .I(N__27662));
    LocalMux I__3787 (
            .O(N__27662),
            .I(\phase_controller_inst1.stoper_tr.counter_i_2 ));
    InMux I__3786 (
            .O(N__27659),
            .I(N__27656));
    LocalMux I__3785 (
            .O(N__27656),
            .I(N__27653));
    Span4Mux_h I__3784 (
            .O(N__27653),
            .I(N__27650));
    Odrv4 I__3783 (
            .O(N__27650),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ));
    InMux I__3782 (
            .O(N__27647),
            .I(N__27643));
    InMux I__3781 (
            .O(N__27646),
            .I(N__27640));
    LocalMux I__3780 (
            .O(N__27643),
            .I(N__27637));
    LocalMux I__3779 (
            .O(N__27640),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ));
    Odrv4 I__3778 (
            .O(N__27637),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ));
    InMux I__3777 (
            .O(N__27632),
            .I(N__27629));
    LocalMux I__3776 (
            .O(N__27629),
            .I(N__27625));
    InMux I__3775 (
            .O(N__27628),
            .I(N__27622));
    Span4Mux_v I__3774 (
            .O(N__27625),
            .I(N__27619));
    LocalMux I__3773 (
            .O(N__27622),
            .I(N__27616));
    Odrv4 I__3772 (
            .O(N__27619),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ));
    Odrv4 I__3771 (
            .O(N__27616),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ));
    InMux I__3770 (
            .O(N__27611),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ));
    InMux I__3769 (
            .O(N__27608),
            .I(N__27605));
    LocalMux I__3768 (
            .O(N__27605),
            .I(N__27602));
    Odrv12 I__3767 (
            .O(N__27602),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ));
    InMux I__3766 (
            .O(N__27599),
            .I(N__27596));
    LocalMux I__3765 (
            .O(N__27596),
            .I(N__27592));
    InMux I__3764 (
            .O(N__27595),
            .I(N__27589));
    Span4Mux_h I__3763 (
            .O(N__27592),
            .I(N__27586));
    LocalMux I__3762 (
            .O(N__27589),
            .I(N__27583));
    Odrv4 I__3761 (
            .O(N__27586),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ));
    Odrv4 I__3760 (
            .O(N__27583),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ));
    InMux I__3759 (
            .O(N__27578),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ));
    InMux I__3758 (
            .O(N__27575),
            .I(N__27571));
    InMux I__3757 (
            .O(N__27574),
            .I(N__27568));
    LocalMux I__3756 (
            .O(N__27571),
            .I(N__27565));
    LocalMux I__3755 (
            .O(N__27568),
            .I(N__27560));
    Span4Mux_h I__3754 (
            .O(N__27565),
            .I(N__27560));
    Odrv4 I__3753 (
            .O(N__27560),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ));
    InMux I__3752 (
            .O(N__27557),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ));
    InMux I__3751 (
            .O(N__27554),
            .I(N__27551));
    LocalMux I__3750 (
            .O(N__27551),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ));
    InMux I__3749 (
            .O(N__27548),
            .I(N__27545));
    LocalMux I__3748 (
            .O(N__27545),
            .I(N__27541));
    InMux I__3747 (
            .O(N__27544),
            .I(N__27538));
    Span4Mux_h I__3746 (
            .O(N__27541),
            .I(N__27533));
    LocalMux I__3745 (
            .O(N__27538),
            .I(N__27533));
    Odrv4 I__3744 (
            .O(N__27533),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ));
    InMux I__3743 (
            .O(N__27530),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ));
    InMux I__3742 (
            .O(N__27527),
            .I(N__27523));
    InMux I__3741 (
            .O(N__27526),
            .I(N__27520));
    LocalMux I__3740 (
            .O(N__27523),
            .I(N__27517));
    LocalMux I__3739 (
            .O(N__27520),
            .I(N__27512));
    Span4Mux_h I__3738 (
            .O(N__27517),
            .I(N__27512));
    Odrv4 I__3737 (
            .O(N__27512),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ));
    InMux I__3736 (
            .O(N__27509),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ));
    InMux I__3735 (
            .O(N__27506),
            .I(N__27502));
    InMux I__3734 (
            .O(N__27505),
            .I(N__27499));
    LocalMux I__3733 (
            .O(N__27502),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ));
    LocalMux I__3732 (
            .O(N__27499),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ));
    InMux I__3731 (
            .O(N__27494),
            .I(bfn_9_17_0_));
    InMux I__3730 (
            .O(N__27491),
            .I(N__27487));
    InMux I__3729 (
            .O(N__27490),
            .I(N__27484));
    LocalMux I__3728 (
            .O(N__27487),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ));
    LocalMux I__3727 (
            .O(N__27484),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ));
    InMux I__3726 (
            .O(N__27479),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ));
    InMux I__3725 (
            .O(N__27476),
            .I(N__27472));
    InMux I__3724 (
            .O(N__27475),
            .I(N__27469));
    LocalMux I__3723 (
            .O(N__27472),
            .I(N__27464));
    LocalMux I__3722 (
            .O(N__27469),
            .I(N__27464));
    Span4Mux_v I__3721 (
            .O(N__27464),
            .I(N__27461));
    Odrv4 I__3720 (
            .O(N__27461),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ));
    InMux I__3719 (
            .O(N__27458),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ));
    InMux I__3718 (
            .O(N__27455),
            .I(N__27452));
    LocalMux I__3717 (
            .O(N__27452),
            .I(N__27448));
    InMux I__3716 (
            .O(N__27451),
            .I(N__27445));
    Span4Mux_v I__3715 (
            .O(N__27448),
            .I(N__27442));
    LocalMux I__3714 (
            .O(N__27445),
            .I(N__27439));
    Odrv4 I__3713 (
            .O(N__27442),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ));
    Odrv4 I__3712 (
            .O(N__27439),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ));
    InMux I__3711 (
            .O(N__27434),
            .I(N__27431));
    LocalMux I__3710 (
            .O(N__27431),
            .I(N__27427));
    InMux I__3709 (
            .O(N__27430),
            .I(N__27424));
    Span4Mux_v I__3708 (
            .O(N__27427),
            .I(N__27421));
    LocalMux I__3707 (
            .O(N__27424),
            .I(N__27418));
    Odrv4 I__3706 (
            .O(N__27421),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ));
    Odrv4 I__3705 (
            .O(N__27418),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ));
    InMux I__3704 (
            .O(N__27413),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ));
    InMux I__3703 (
            .O(N__27410),
            .I(N__27407));
    LocalMux I__3702 (
            .O(N__27407),
            .I(N__27403));
    InMux I__3701 (
            .O(N__27406),
            .I(N__27400));
    Span4Mux_h I__3700 (
            .O(N__27403),
            .I(N__27397));
    LocalMux I__3699 (
            .O(N__27400),
            .I(N__27394));
    Odrv4 I__3698 (
            .O(N__27397),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ));
    Odrv4 I__3697 (
            .O(N__27394),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ));
    InMux I__3696 (
            .O(N__27389),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ));
    InMux I__3695 (
            .O(N__27386),
            .I(N__27383));
    LocalMux I__3694 (
            .O(N__27383),
            .I(N__27380));
    Span4Mux_v I__3693 (
            .O(N__27380),
            .I(N__27377));
    Odrv4 I__3692 (
            .O(N__27377),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ));
    InMux I__3691 (
            .O(N__27374),
            .I(N__27370));
    InMux I__3690 (
            .O(N__27373),
            .I(N__27367));
    LocalMux I__3689 (
            .O(N__27370),
            .I(N__27364));
    LocalMux I__3688 (
            .O(N__27367),
            .I(N__27359));
    Span4Mux_h I__3687 (
            .O(N__27364),
            .I(N__27359));
    Odrv4 I__3686 (
            .O(N__27359),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ));
    InMux I__3685 (
            .O(N__27356),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ));
    CascadeMux I__3684 (
            .O(N__27353),
            .I(N__27350));
    InMux I__3683 (
            .O(N__27350),
            .I(N__27347));
    LocalMux I__3682 (
            .O(N__27347),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ));
    InMux I__3681 (
            .O(N__27344),
            .I(N__27341));
    LocalMux I__3680 (
            .O(N__27341),
            .I(N__27337));
    InMux I__3679 (
            .O(N__27340),
            .I(N__27334));
    Span4Mux_h I__3678 (
            .O(N__27337),
            .I(N__27331));
    LocalMux I__3677 (
            .O(N__27334),
            .I(N__27328));
    Odrv4 I__3676 (
            .O(N__27331),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ));
    Odrv4 I__3675 (
            .O(N__27328),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ));
    InMux I__3674 (
            .O(N__27323),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ));
    InMux I__3673 (
            .O(N__27320),
            .I(N__27316));
    InMux I__3672 (
            .O(N__27319),
            .I(N__27313));
    LocalMux I__3671 (
            .O(N__27316),
            .I(N__27310));
    LocalMux I__3670 (
            .O(N__27313),
            .I(N__27305));
    Span4Mux_h I__3669 (
            .O(N__27310),
            .I(N__27305));
    Odrv4 I__3668 (
            .O(N__27305),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ));
    InMux I__3667 (
            .O(N__27302),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ));
    InMux I__3666 (
            .O(N__27299),
            .I(N__27295));
    InMux I__3665 (
            .O(N__27298),
            .I(N__27292));
    LocalMux I__3664 (
            .O(N__27295),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ));
    LocalMux I__3663 (
            .O(N__27292),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ));
    InMux I__3662 (
            .O(N__27287),
            .I(bfn_9_16_0_));
    InMux I__3661 (
            .O(N__27284),
            .I(N__27280));
    InMux I__3660 (
            .O(N__27283),
            .I(N__27277));
    LocalMux I__3659 (
            .O(N__27280),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ));
    LocalMux I__3658 (
            .O(N__27277),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ));
    InMux I__3657 (
            .O(N__27272),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ));
    InMux I__3656 (
            .O(N__27269),
            .I(N__27265));
    InMux I__3655 (
            .O(N__27268),
            .I(N__27262));
    LocalMux I__3654 (
            .O(N__27265),
            .I(N__27259));
    LocalMux I__3653 (
            .O(N__27262),
            .I(N__27256));
    Span4Mux_v I__3652 (
            .O(N__27259),
            .I(N__27253));
    Odrv4 I__3651 (
            .O(N__27256),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ));
    Odrv4 I__3650 (
            .O(N__27253),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ));
    InMux I__3649 (
            .O(N__27248),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ));
    InMux I__3648 (
            .O(N__27245),
            .I(N__27242));
    LocalMux I__3647 (
            .O(N__27242),
            .I(N__27238));
    InMux I__3646 (
            .O(N__27241),
            .I(N__27235));
    Span4Mux_v I__3645 (
            .O(N__27238),
            .I(N__27232));
    LocalMux I__3644 (
            .O(N__27235),
            .I(N__27229));
    Odrv4 I__3643 (
            .O(N__27232),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ));
    Odrv4 I__3642 (
            .O(N__27229),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ));
    InMux I__3641 (
            .O(N__27224),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ));
    InMux I__3640 (
            .O(N__27221),
            .I(N__27217));
    InMux I__3639 (
            .O(N__27220),
            .I(N__27214));
    LocalMux I__3638 (
            .O(N__27217),
            .I(N__27209));
    LocalMux I__3637 (
            .O(N__27214),
            .I(N__27209));
    Span4Mux_h I__3636 (
            .O(N__27209),
            .I(N__27206));
    Odrv4 I__3635 (
            .O(N__27206),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ));
    InMux I__3634 (
            .O(N__27203),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ));
    InMux I__3633 (
            .O(N__27200),
            .I(N__27196));
    InMux I__3632 (
            .O(N__27199),
            .I(N__27193));
    LocalMux I__3631 (
            .O(N__27196),
            .I(N__27190));
    LocalMux I__3630 (
            .O(N__27193),
            .I(N__27185));
    Span4Mux_h I__3629 (
            .O(N__27190),
            .I(N__27185));
    Odrv4 I__3628 (
            .O(N__27185),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ));
    InMux I__3627 (
            .O(N__27182),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ));
    InMux I__3626 (
            .O(N__27179),
            .I(N__27176));
    LocalMux I__3625 (
            .O(N__27176),
            .I(N__27173));
    Odrv4 I__3624 (
            .O(N__27173),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ));
    InMux I__3623 (
            .O(N__27170),
            .I(N__27167));
    LocalMux I__3622 (
            .O(N__27167),
            .I(N__27163));
    InMux I__3621 (
            .O(N__27166),
            .I(N__27160));
    Span4Mux_h I__3620 (
            .O(N__27163),
            .I(N__27157));
    LocalMux I__3619 (
            .O(N__27160),
            .I(N__27154));
    Odrv4 I__3618 (
            .O(N__27157),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ));
    Odrv4 I__3617 (
            .O(N__27154),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ));
    InMux I__3616 (
            .O(N__27149),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ));
    InMux I__3615 (
            .O(N__27146),
            .I(N__27142));
    InMux I__3614 (
            .O(N__27145),
            .I(N__27139));
    LocalMux I__3613 (
            .O(N__27142),
            .I(N__27136));
    LocalMux I__3612 (
            .O(N__27139),
            .I(N__27131));
    Span4Mux_h I__3611 (
            .O(N__27136),
            .I(N__27131));
    Odrv4 I__3610 (
            .O(N__27131),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ));
    InMux I__3609 (
            .O(N__27128),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ));
    InMux I__3608 (
            .O(N__27125),
            .I(N__27121));
    InMux I__3607 (
            .O(N__27124),
            .I(N__27118));
    LocalMux I__3606 (
            .O(N__27121),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ));
    LocalMux I__3605 (
            .O(N__27118),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ));
    InMux I__3604 (
            .O(N__27113),
            .I(bfn_9_15_0_));
    InMux I__3603 (
            .O(N__27110),
            .I(N__27106));
    InMux I__3602 (
            .O(N__27109),
            .I(N__27103));
    LocalMux I__3601 (
            .O(N__27106),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ));
    LocalMux I__3600 (
            .O(N__27103),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ));
    InMux I__3599 (
            .O(N__27098),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ));
    InMux I__3598 (
            .O(N__27095),
            .I(N__27091));
    InMux I__3597 (
            .O(N__27094),
            .I(N__27088));
    LocalMux I__3596 (
            .O(N__27091),
            .I(N__27083));
    LocalMux I__3595 (
            .O(N__27088),
            .I(N__27083));
    Span4Mux_v I__3594 (
            .O(N__27083),
            .I(N__27080));
    Odrv4 I__3593 (
            .O(N__27080),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ));
    InMux I__3592 (
            .O(N__27077),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ));
    InMux I__3591 (
            .O(N__27074),
            .I(N__27068));
    InMux I__3590 (
            .O(N__27073),
            .I(N__27068));
    LocalMux I__3589 (
            .O(N__27068),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__3588 (
            .O(N__27065),
            .I(N__27059));
    InMux I__3587 (
            .O(N__27064),
            .I(N__27059));
    LocalMux I__3586 (
            .O(N__27059),
            .I(N__27056));
    Odrv4 I__3585 (
            .O(N__27056),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__3584 (
            .O(N__27053),
            .I(N__27050));
    LocalMux I__3583 (
            .O(N__27050),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    CascadeMux I__3582 (
            .O(N__27047),
            .I(elapsed_time_ns_1_RNIFE91B_0_3_cascade_));
    InMux I__3581 (
            .O(N__27044),
            .I(N__27040));
    InMux I__3580 (
            .O(N__27043),
            .I(N__27037));
    LocalMux I__3579 (
            .O(N__27040),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__3578 (
            .O(N__27037),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    CascadeMux I__3577 (
            .O(N__27032),
            .I(N__27029));
    InMux I__3576 (
            .O(N__27029),
            .I(N__27026));
    LocalMux I__3575 (
            .O(N__27026),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ));
    InMux I__3574 (
            .O(N__27023),
            .I(N__27019));
    InMux I__3573 (
            .O(N__27022),
            .I(N__27016));
    LocalMux I__3572 (
            .O(N__27019),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    LocalMux I__3571 (
            .O(N__27016),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__3570 (
            .O(N__27011),
            .I(N__27008));
    LocalMux I__3569 (
            .O(N__27008),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ));
    InMux I__3568 (
            .O(N__27005),
            .I(N__27002));
    LocalMux I__3567 (
            .O(N__27002),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ));
    InMux I__3566 (
            .O(N__26999),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ));
    InMux I__3565 (
            .O(N__26996),
            .I(N__26993));
    LocalMux I__3564 (
            .O(N__26993),
            .I(N__26989));
    InMux I__3563 (
            .O(N__26992),
            .I(N__26986));
    Span4Mux_s1_v I__3562 (
            .O(N__26989),
            .I(N__26981));
    LocalMux I__3561 (
            .O(N__26986),
            .I(N__26981));
    Span4Mux_v I__3560 (
            .O(N__26981),
            .I(N__26977));
    InMux I__3559 (
            .O(N__26980),
            .I(N__26972));
    Span4Mux_h I__3558 (
            .O(N__26977),
            .I(N__26966));
    InMux I__3557 (
            .O(N__26976),
            .I(N__26961));
    InMux I__3556 (
            .O(N__26975),
            .I(N__26961));
    LocalMux I__3555 (
            .O(N__26972),
            .I(N__26958));
    InMux I__3554 (
            .O(N__26971),
            .I(N__26951));
    InMux I__3553 (
            .O(N__26970),
            .I(N__26951));
    InMux I__3552 (
            .O(N__26969),
            .I(N__26951));
    Sp12to4 I__3551 (
            .O(N__26966),
            .I(N__26948));
    LocalMux I__3550 (
            .O(N__26961),
            .I(N__26945));
    Span4Mux_v I__3549 (
            .O(N__26958),
            .I(N__26940));
    LocalMux I__3548 (
            .O(N__26951),
            .I(N__26940));
    Span12Mux_s11_v I__3547 (
            .O(N__26948),
            .I(N__26937));
    Span4Mux_v I__3546 (
            .O(N__26945),
            .I(N__26934));
    Span4Mux_v I__3545 (
            .O(N__26940),
            .I(N__26931));
    Span12Mux_v I__3544 (
            .O(N__26937),
            .I(N__26924));
    Sp12to4 I__3543 (
            .O(N__26934),
            .I(N__26924));
    Sp12to4 I__3542 (
            .O(N__26931),
            .I(N__26924));
    Span12Mux_h I__3541 (
            .O(N__26924),
            .I(N__26921));
    Odrv12 I__3540 (
            .O(N__26921),
            .I(start_stop_c));
    InMux I__3539 (
            .O(N__26918),
            .I(N__26914));
    CascadeMux I__3538 (
            .O(N__26917),
            .I(N__26911));
    LocalMux I__3537 (
            .O(N__26914),
            .I(N__26907));
    InMux I__3536 (
            .O(N__26911),
            .I(N__26902));
    InMux I__3535 (
            .O(N__26910),
            .I(N__26902));
    Span4Mux_h I__3534 (
            .O(N__26907),
            .I(N__26899));
    LocalMux I__3533 (
            .O(N__26902),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    Odrv4 I__3532 (
            .O(N__26899),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    CascadeMux I__3531 (
            .O(N__26894),
            .I(\phase_controller_inst1.state_ns_0_0_1_cascade_ ));
    InMux I__3530 (
            .O(N__26891),
            .I(N__26888));
    LocalMux I__3529 (
            .O(N__26888),
            .I(N__26885));
    Span4Mux_h I__3528 (
            .O(N__26885),
            .I(N__26880));
    InMux I__3527 (
            .O(N__26884),
            .I(N__26875));
    InMux I__3526 (
            .O(N__26883),
            .I(N__26875));
    Odrv4 I__3525 (
            .O(N__26880),
            .I(\phase_controller_inst1.start_flagZ0 ));
    LocalMux I__3524 (
            .O(N__26875),
            .I(\phase_controller_inst1.start_flagZ0 ));
    CascadeMux I__3523 (
            .O(N__26870),
            .I(\phase_controller_inst1.stoper_tr.un4_start_0_cascade_ ));
    CascadeMux I__3522 (
            .O(N__26867),
            .I(N__26862));
    InMux I__3521 (
            .O(N__26866),
            .I(N__26855));
    InMux I__3520 (
            .O(N__26865),
            .I(N__26855));
    InMux I__3519 (
            .O(N__26862),
            .I(N__26855));
    LocalMux I__3518 (
            .O(N__26855),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__3517 (
            .O(N__26852),
            .I(N__26846));
    InMux I__3516 (
            .O(N__26851),
            .I(N__26846));
    LocalMux I__3515 (
            .O(N__26846),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__3514 (
            .O(N__26843),
            .I(N__26840));
    LocalMux I__3513 (
            .O(N__26840),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    CascadeMux I__3512 (
            .O(N__26837),
            .I(elapsed_time_ns_1_RNIJI91B_0_7_cascade_));
    InMux I__3511 (
            .O(N__26834),
            .I(N__26830));
    InMux I__3510 (
            .O(N__26833),
            .I(N__26827));
    LocalMux I__3509 (
            .O(N__26830),
            .I(N__26824));
    LocalMux I__3508 (
            .O(N__26827),
            .I(N__26821));
    Span4Mux_h I__3507 (
            .O(N__26824),
            .I(N__26817));
    Span4Mux_h I__3506 (
            .O(N__26821),
            .I(N__26814));
    InMux I__3505 (
            .O(N__26820),
            .I(N__26811));
    Span4Mux_v I__3504 (
            .O(N__26817),
            .I(N__26808));
    Sp12to4 I__3503 (
            .O(N__26814),
            .I(N__26803));
    LocalMux I__3502 (
            .O(N__26811),
            .I(N__26803));
    Odrv4 I__3501 (
            .O(N__26808),
            .I(il_min_comp2_c));
    Odrv12 I__3500 (
            .O(N__26803),
            .I(il_min_comp2_c));
    InMux I__3499 (
            .O(N__26798),
            .I(N__26794));
    CascadeMux I__3498 (
            .O(N__26797),
            .I(N__26791));
    LocalMux I__3497 (
            .O(N__26794),
            .I(N__26788));
    InMux I__3496 (
            .O(N__26791),
            .I(N__26783));
    Sp12to4 I__3495 (
            .O(N__26788),
            .I(N__26780));
    InMux I__3494 (
            .O(N__26787),
            .I(N__26777));
    InMux I__3493 (
            .O(N__26786),
            .I(N__26774));
    LocalMux I__3492 (
            .O(N__26783),
            .I(N__26771));
    Span12Mux_v I__3491 (
            .O(N__26780),
            .I(N__26768));
    LocalMux I__3490 (
            .O(N__26777),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__3489 (
            .O(N__26774),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__3488 (
            .O(N__26771),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv12 I__3487 (
            .O(N__26768),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__3486 (
            .O(N__26759),
            .I(N__26753));
    InMux I__3485 (
            .O(N__26758),
            .I(N__26753));
    LocalMux I__3484 (
            .O(N__26753),
            .I(N__26749));
    InMux I__3483 (
            .O(N__26752),
            .I(N__26746));
    Span4Mux_v I__3482 (
            .O(N__26749),
            .I(N__26741));
    LocalMux I__3481 (
            .O(N__26746),
            .I(N__26741));
    Span4Mux_v I__3480 (
            .O(N__26741),
            .I(N__26738));
    Span4Mux_h I__3479 (
            .O(N__26738),
            .I(N__26735));
    Odrv4 I__3478 (
            .O(N__26735),
            .I(il_max_comp2_c));
    CascadeMux I__3477 (
            .O(N__26732),
            .I(N__26727));
    CascadeMux I__3476 (
            .O(N__26731),
            .I(N__26724));
    InMux I__3475 (
            .O(N__26730),
            .I(N__26716));
    InMux I__3474 (
            .O(N__26727),
            .I(N__26716));
    InMux I__3473 (
            .O(N__26724),
            .I(N__26716));
    InMux I__3472 (
            .O(N__26723),
            .I(N__26713));
    LocalMux I__3471 (
            .O(N__26716),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__3470 (
            .O(N__26713),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__3469 (
            .O(N__26708),
            .I(N__26699));
    InMux I__3468 (
            .O(N__26707),
            .I(N__26699));
    InMux I__3467 (
            .O(N__26706),
            .I(N__26691));
    InMux I__3466 (
            .O(N__26705),
            .I(N__26691));
    InMux I__3465 (
            .O(N__26704),
            .I(N__26691));
    LocalMux I__3464 (
            .O(N__26699),
            .I(N__26688));
    InMux I__3463 (
            .O(N__26698),
            .I(N__26685));
    LocalMux I__3462 (
            .O(N__26691),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__3461 (
            .O(N__26688),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__3460 (
            .O(N__26685),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__3459 (
            .O(N__26678),
            .I(N__26673));
    InMux I__3458 (
            .O(N__26677),
            .I(N__26668));
    InMux I__3457 (
            .O(N__26676),
            .I(N__26668));
    LocalMux I__3456 (
            .O(N__26673),
            .I(N__26665));
    LocalMux I__3455 (
            .O(N__26668),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    Odrv4 I__3454 (
            .O(N__26665),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__3453 (
            .O(N__26660),
            .I(N__26657));
    LocalMux I__3452 (
            .O(N__26657),
            .I(\phase_controller_inst2.stoper_hc.un4_start_0 ));
    InMux I__3451 (
            .O(N__26654),
            .I(N__26644));
    InMux I__3450 (
            .O(N__26653),
            .I(N__26644));
    InMux I__3449 (
            .O(N__26652),
            .I(N__26644));
    InMux I__3448 (
            .O(N__26651),
            .I(N__26641));
    LocalMux I__3447 (
            .O(N__26644),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__3446 (
            .O(N__26641),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__3445 (
            .O(N__26636),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_28 ));
    InMux I__3444 (
            .O(N__26633),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_29 ));
    InMux I__3443 (
            .O(N__26630),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_30 ));
    CEMux I__3442 (
            .O(N__26627),
            .I(N__26615));
    CEMux I__3441 (
            .O(N__26626),
            .I(N__26615));
    CEMux I__3440 (
            .O(N__26625),
            .I(N__26615));
    CEMux I__3439 (
            .O(N__26624),
            .I(N__26615));
    GlobalMux I__3438 (
            .O(N__26615),
            .I(N__26612));
    gio2CtrlBuf I__3437 (
            .O(N__26612),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0_g ));
    IoInMux I__3436 (
            .O(N__26609),
            .I(N__26606));
    LocalMux I__3435 (
            .O(N__26606),
            .I(N__26603));
    Odrv12 I__3434 (
            .O(N__26603),
            .I(s4_phy_c));
    CascadeMux I__3433 (
            .O(N__26600),
            .I(N__26596));
    CascadeMux I__3432 (
            .O(N__26599),
            .I(N__26592));
    InMux I__3431 (
            .O(N__26596),
            .I(N__26589));
    InMux I__3430 (
            .O(N__26595),
            .I(N__26586));
    InMux I__3429 (
            .O(N__26592),
            .I(N__26583));
    LocalMux I__3428 (
            .O(N__26589),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__3427 (
            .O(N__26586),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__3426 (
            .O(N__26583),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__3425 (
            .O(N__26576),
            .I(N__26572));
    InMux I__3424 (
            .O(N__26575),
            .I(N__26569));
    LocalMux I__3423 (
            .O(N__26572),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__3422 (
            .O(N__26569),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__3421 (
            .O(N__26564),
            .I(N__26561));
    LocalMux I__3420 (
            .O(N__26561),
            .I(\phase_controller_inst2.state_ns_0_0_1 ));
    InMux I__3419 (
            .O(N__26558),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_19 ));
    InMux I__3418 (
            .O(N__26555),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_20 ));
    InMux I__3417 (
            .O(N__26552),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_21 ));
    InMux I__3416 (
            .O(N__26549),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_22 ));
    InMux I__3415 (
            .O(N__26546),
            .I(bfn_8_23_0_));
    InMux I__3414 (
            .O(N__26543),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_24 ));
    InMux I__3413 (
            .O(N__26540),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_25 ));
    InMux I__3412 (
            .O(N__26537),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_26 ));
    InMux I__3411 (
            .O(N__26534),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_27 ));
    InMux I__3410 (
            .O(N__26531),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_10 ));
    InMux I__3409 (
            .O(N__26528),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_11 ));
    InMux I__3408 (
            .O(N__26525),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_12 ));
    InMux I__3407 (
            .O(N__26522),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_13 ));
    InMux I__3406 (
            .O(N__26519),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_14 ));
    InMux I__3405 (
            .O(N__26516),
            .I(bfn_8_22_0_));
    InMux I__3404 (
            .O(N__26513),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_16 ));
    CascadeMux I__3403 (
            .O(N__26510),
            .I(N__26506));
    CascadeMux I__3402 (
            .O(N__26509),
            .I(N__26503));
    InMux I__3401 (
            .O(N__26506),
            .I(N__26497));
    InMux I__3400 (
            .O(N__26503),
            .I(N__26497));
    InMux I__3399 (
            .O(N__26502),
            .I(N__26494));
    LocalMux I__3398 (
            .O(N__26497),
            .I(N__26491));
    LocalMux I__3397 (
            .O(N__26494),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ));
    Odrv4 I__3396 (
            .O(N__26491),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ));
    InMux I__3395 (
            .O(N__26486),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_17 ));
    InMux I__3394 (
            .O(N__26483),
            .I(N__26476));
    InMux I__3393 (
            .O(N__26482),
            .I(N__26476));
    InMux I__3392 (
            .O(N__26481),
            .I(N__26473));
    LocalMux I__3391 (
            .O(N__26476),
            .I(N__26470));
    LocalMux I__3390 (
            .O(N__26473),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ));
    Odrv4 I__3389 (
            .O(N__26470),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ));
    InMux I__3388 (
            .O(N__26465),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_18 ));
    InMux I__3387 (
            .O(N__26462),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_1 ));
    InMux I__3386 (
            .O(N__26459),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_2 ));
    InMux I__3385 (
            .O(N__26456),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_3 ));
    InMux I__3384 (
            .O(N__26453),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_4 ));
    InMux I__3383 (
            .O(N__26450),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_5 ));
    InMux I__3382 (
            .O(N__26447),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_6 ));
    InMux I__3381 (
            .O(N__26444),
            .I(bfn_8_21_0_));
    InMux I__3380 (
            .O(N__26441),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_8 ));
    InMux I__3379 (
            .O(N__26438),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_9 ));
    InMux I__3378 (
            .O(N__26435),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ));
    InMux I__3377 (
            .O(N__26432),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ));
    InMux I__3376 (
            .O(N__26429),
            .I(bfn_8_19_0_));
    InMux I__3375 (
            .O(N__26426),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ));
    InMux I__3374 (
            .O(N__26423),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ));
    InMux I__3373 (
            .O(N__26420),
            .I(N__26417));
    LocalMux I__3372 (
            .O(N__26417),
            .I(N__26413));
    InMux I__3371 (
            .O(N__26416),
            .I(N__26410));
    Span4Mux_v I__3370 (
            .O(N__26413),
            .I(N__26405));
    LocalMux I__3369 (
            .O(N__26410),
            .I(N__26405));
    Odrv4 I__3368 (
            .O(N__26405),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_27));
    InMux I__3367 (
            .O(N__26402),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ));
    InMux I__3366 (
            .O(N__26399),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ));
    InMux I__3365 (
            .O(N__26396),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_0 ));
    InMux I__3364 (
            .O(N__26393),
            .I(N__26390));
    LocalMux I__3363 (
            .O(N__26390),
            .I(N__26387));
    Span4Mux_h I__3362 (
            .O(N__26387),
            .I(N__26383));
    InMux I__3361 (
            .O(N__26386),
            .I(N__26380));
    Odrv4 I__3360 (
            .O(N__26383),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_13));
    LocalMux I__3359 (
            .O(N__26380),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_13));
    InMux I__3358 (
            .O(N__26375),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ));
    InMux I__3357 (
            .O(N__26372),
            .I(N__26369));
    LocalMux I__3356 (
            .O(N__26369),
            .I(N__26366));
    Span4Mux_h I__3355 (
            .O(N__26366),
            .I(N__26362));
    InMux I__3354 (
            .O(N__26365),
            .I(N__26359));
    Odrv4 I__3353 (
            .O(N__26362),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_14));
    LocalMux I__3352 (
            .O(N__26359),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_14));
    InMux I__3351 (
            .O(N__26354),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ));
    InMux I__3350 (
            .O(N__26351),
            .I(N__26348));
    LocalMux I__3349 (
            .O(N__26348),
            .I(N__26345));
    Span4Mux_v I__3348 (
            .O(N__26345),
            .I(N__26341));
    InMux I__3347 (
            .O(N__26344),
            .I(N__26338));
    Odrv4 I__3346 (
            .O(N__26341),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_15));
    LocalMux I__3345 (
            .O(N__26338),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_15));
    InMux I__3344 (
            .O(N__26333),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ));
    InMux I__3343 (
            .O(N__26330),
            .I(N__26326));
    InMux I__3342 (
            .O(N__26329),
            .I(N__26323));
    LocalMux I__3341 (
            .O(N__26326),
            .I(N__26320));
    LocalMux I__3340 (
            .O(N__26323),
            .I(N__26317));
    Odrv4 I__3339 (
            .O(N__26320),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_16));
    Odrv4 I__3338 (
            .O(N__26317),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_16));
    InMux I__3337 (
            .O(N__26312),
            .I(bfn_8_18_0_));
    InMux I__3336 (
            .O(N__26309),
            .I(N__26305));
    InMux I__3335 (
            .O(N__26308),
            .I(N__26302));
    LocalMux I__3334 (
            .O(N__26305),
            .I(N__26299));
    LocalMux I__3333 (
            .O(N__26302),
            .I(N__26296));
    Odrv4 I__3332 (
            .O(N__26299),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_17));
    Odrv4 I__3331 (
            .O(N__26296),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_17));
    InMux I__3330 (
            .O(N__26291),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ));
    InMux I__3329 (
            .O(N__26288),
            .I(N__26285));
    LocalMux I__3328 (
            .O(N__26285),
            .I(N__26281));
    InMux I__3327 (
            .O(N__26284),
            .I(N__26278));
    Span4Mux_v I__3326 (
            .O(N__26281),
            .I(N__26273));
    LocalMux I__3325 (
            .O(N__26278),
            .I(N__26273));
    Odrv4 I__3324 (
            .O(N__26273),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_18));
    InMux I__3323 (
            .O(N__26270),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ));
    InMux I__3322 (
            .O(N__26267),
            .I(N__26264));
    LocalMux I__3321 (
            .O(N__26264),
            .I(N__26260));
    InMux I__3320 (
            .O(N__26263),
            .I(N__26257));
    Span4Mux_v I__3319 (
            .O(N__26260),
            .I(N__26252));
    LocalMux I__3318 (
            .O(N__26257),
            .I(N__26252));
    Odrv4 I__3317 (
            .O(N__26252),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_19));
    InMux I__3316 (
            .O(N__26249),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ));
    InMux I__3315 (
            .O(N__26246),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ));
    InMux I__3314 (
            .O(N__26243),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ));
    InMux I__3313 (
            .O(N__26240),
            .I(N__26237));
    LocalMux I__3312 (
            .O(N__26237),
            .I(N__26233));
    InMux I__3311 (
            .O(N__26236),
            .I(N__26230));
    Odrv4 I__3310 (
            .O(N__26233),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_5));
    LocalMux I__3309 (
            .O(N__26230),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_5));
    InMux I__3308 (
            .O(N__26225),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ));
    InMux I__3307 (
            .O(N__26222),
            .I(N__26219));
    LocalMux I__3306 (
            .O(N__26219),
            .I(N__26215));
    InMux I__3305 (
            .O(N__26218),
            .I(N__26212));
    Odrv4 I__3304 (
            .O(N__26215),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_6));
    LocalMux I__3303 (
            .O(N__26212),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_6));
    InMux I__3302 (
            .O(N__26207),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ));
    InMux I__3301 (
            .O(N__26204),
            .I(N__26200));
    InMux I__3300 (
            .O(N__26203),
            .I(N__26197));
    LocalMux I__3299 (
            .O(N__26200),
            .I(N__26194));
    LocalMux I__3298 (
            .O(N__26197),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_7));
    Odrv4 I__3297 (
            .O(N__26194),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_7));
    InMux I__3296 (
            .O(N__26189),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ));
    InMux I__3295 (
            .O(N__26186),
            .I(N__26182));
    InMux I__3294 (
            .O(N__26185),
            .I(N__26179));
    LocalMux I__3293 (
            .O(N__26182),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_8));
    LocalMux I__3292 (
            .O(N__26179),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_8));
    InMux I__3291 (
            .O(N__26174),
            .I(bfn_8_17_0_));
    InMux I__3290 (
            .O(N__26171),
            .I(N__26168));
    LocalMux I__3289 (
            .O(N__26168),
            .I(N__26164));
    InMux I__3288 (
            .O(N__26167),
            .I(N__26161));
    Odrv4 I__3287 (
            .O(N__26164),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_9));
    LocalMux I__3286 (
            .O(N__26161),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_9));
    InMux I__3285 (
            .O(N__26156),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ));
    InMux I__3284 (
            .O(N__26153),
            .I(N__26149));
    InMux I__3283 (
            .O(N__26152),
            .I(N__26146));
    LocalMux I__3282 (
            .O(N__26149),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_10));
    LocalMux I__3281 (
            .O(N__26146),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_10));
    InMux I__3280 (
            .O(N__26141),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ));
    InMux I__3279 (
            .O(N__26138),
            .I(N__26135));
    LocalMux I__3278 (
            .O(N__26135),
            .I(N__26131));
    InMux I__3277 (
            .O(N__26134),
            .I(N__26128));
    Odrv4 I__3276 (
            .O(N__26131),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_11));
    LocalMux I__3275 (
            .O(N__26128),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_11));
    InMux I__3274 (
            .O(N__26123),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ));
    InMux I__3273 (
            .O(N__26120),
            .I(N__26117));
    LocalMux I__3272 (
            .O(N__26117),
            .I(N__26114));
    Span4Mux_h I__3271 (
            .O(N__26114),
            .I(N__26110));
    InMux I__3270 (
            .O(N__26113),
            .I(N__26107));
    Odrv4 I__3269 (
            .O(N__26110),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_12));
    LocalMux I__3268 (
            .O(N__26107),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_12));
    InMux I__3267 (
            .O(N__26102),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ));
    InMux I__3266 (
            .O(N__26099),
            .I(N__26096));
    LocalMux I__3265 (
            .O(N__26096),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    CascadeMux I__3264 (
            .O(N__26093),
            .I(elapsed_time_ns_1_RNI2COBB_0_15_cascade_));
    InMux I__3263 (
            .O(N__26090),
            .I(N__26086));
    InMux I__3262 (
            .O(N__26089),
            .I(N__26083));
    LocalMux I__3261 (
            .O(N__26086),
            .I(N__26080));
    LocalMux I__3260 (
            .O(N__26083),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    Odrv4 I__3259 (
            .O(N__26080),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    CascadeMux I__3258 (
            .O(N__26075),
            .I(N__26072));
    InMux I__3257 (
            .O(N__26072),
            .I(N__26069));
    LocalMux I__3256 (
            .O(N__26069),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt30 ));
    InMux I__3255 (
            .O(N__26066),
            .I(N__26063));
    LocalMux I__3254 (
            .O(N__26063),
            .I(\phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ));
    InMux I__3253 (
            .O(N__26060),
            .I(N__26056));
    InMux I__3252 (
            .O(N__26059),
            .I(N__26053));
    LocalMux I__3251 (
            .O(N__26056),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_1));
    LocalMux I__3250 (
            .O(N__26053),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_1));
    InMux I__3249 (
            .O(N__26048),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ));
    InMux I__3248 (
            .O(N__26045),
            .I(N__26042));
    LocalMux I__3247 (
            .O(N__26042),
            .I(N__26038));
    InMux I__3246 (
            .O(N__26041),
            .I(N__26035));
    Odrv4 I__3245 (
            .O(N__26038),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_2));
    LocalMux I__3244 (
            .O(N__26035),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_2));
    InMux I__3243 (
            .O(N__26030),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ));
    InMux I__3242 (
            .O(N__26027),
            .I(N__26023));
    InMux I__3241 (
            .O(N__26026),
            .I(N__26020));
    LocalMux I__3240 (
            .O(N__26023),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_3));
    LocalMux I__3239 (
            .O(N__26020),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_3));
    InMux I__3238 (
            .O(N__26015),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ));
    InMux I__3237 (
            .O(N__26012),
            .I(N__26009));
    LocalMux I__3236 (
            .O(N__26009),
            .I(N__26005));
    InMux I__3235 (
            .O(N__26008),
            .I(N__26002));
    Odrv4 I__3234 (
            .O(N__26005),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_4));
    LocalMux I__3233 (
            .O(N__26002),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_4));
    InMux I__3232 (
            .O(N__25997),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ));
    InMux I__3231 (
            .O(N__25994),
            .I(N__25991));
    LocalMux I__3230 (
            .O(N__25991),
            .I(N__25988));
    Odrv4 I__3229 (
            .O(N__25988),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ));
    CascadeMux I__3228 (
            .O(N__25985),
            .I(N__25982));
    InMux I__3227 (
            .O(N__25982),
            .I(N__25979));
    LocalMux I__3226 (
            .O(N__25979),
            .I(N__25976));
    Span4Mux_h I__3225 (
            .O(N__25976),
            .I(N__25973));
    Odrv4 I__3224 (
            .O(N__25973),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt24 ));
    InMux I__3223 (
            .O(N__25970),
            .I(N__25967));
    LocalMux I__3222 (
            .O(N__25967),
            .I(N__25964));
    Odrv4 I__3221 (
            .O(N__25964),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt26 ));
    CascadeMux I__3220 (
            .O(N__25961),
            .I(N__25958));
    InMux I__3219 (
            .O(N__25958),
            .I(N__25955));
    LocalMux I__3218 (
            .O(N__25955),
            .I(N__25952));
    Span4Mux_v I__3217 (
            .O(N__25952),
            .I(N__25949));
    Odrv4 I__3216 (
            .O(N__25949),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ));
    InMux I__3215 (
            .O(N__25946),
            .I(bfn_8_15_0_));
    CascadeMux I__3214 (
            .O(N__25943),
            .I(N__25940));
    InMux I__3213 (
            .O(N__25940),
            .I(N__25937));
    LocalMux I__3212 (
            .O(N__25937),
            .I(N__25934));
    Odrv4 I__3211 (
            .O(N__25934),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt28 ));
    InMux I__3210 (
            .O(N__25931),
            .I(N__25925));
    InMux I__3209 (
            .O(N__25930),
            .I(N__25925));
    LocalMux I__3208 (
            .O(N__25925),
            .I(N__25921));
    InMux I__3207 (
            .O(N__25924),
            .I(N__25918));
    Span4Mux_v I__3206 (
            .O(N__25921),
            .I(N__25915));
    LocalMux I__3205 (
            .O(N__25918),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ));
    Odrv4 I__3204 (
            .O(N__25915),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ));
    CascadeMux I__3203 (
            .O(N__25910),
            .I(N__25907));
    InMux I__3202 (
            .O(N__25907),
            .I(N__25901));
    InMux I__3201 (
            .O(N__25906),
            .I(N__25901));
    LocalMux I__3200 (
            .O(N__25901),
            .I(N__25897));
    InMux I__3199 (
            .O(N__25900),
            .I(N__25894));
    Span4Mux_v I__3198 (
            .O(N__25897),
            .I(N__25891));
    LocalMux I__3197 (
            .O(N__25894),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ));
    Odrv4 I__3196 (
            .O(N__25891),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ));
    InMux I__3195 (
            .O(N__25886),
            .I(N__25883));
    LocalMux I__3194 (
            .O(N__25883),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ));
    InMux I__3193 (
            .O(N__25880),
            .I(N__25877));
    LocalMux I__3192 (
            .O(N__25877),
            .I(N__25870));
    CascadeMux I__3191 (
            .O(N__25876),
            .I(N__25867));
    InMux I__3190 (
            .O(N__25875),
            .I(N__25861));
    InMux I__3189 (
            .O(N__25874),
            .I(N__25861));
    InMux I__3188 (
            .O(N__25873),
            .I(N__25858));
    Span4Mux_v I__3187 (
            .O(N__25870),
            .I(N__25855));
    InMux I__3186 (
            .O(N__25867),
            .I(N__25852));
    InMux I__3185 (
            .O(N__25866),
            .I(N__25849));
    LocalMux I__3184 (
            .O(N__25861),
            .I(N__25846));
    LocalMux I__3183 (
            .O(N__25858),
            .I(N__25843));
    Span4Mux_v I__3182 (
            .O(N__25855),
            .I(N__25840));
    LocalMux I__3181 (
            .O(N__25852),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__3180 (
            .O(N__25849),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__3179 (
            .O(N__25846),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__3178 (
            .O(N__25843),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__3177 (
            .O(N__25840),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__3176 (
            .O(N__25829),
            .I(N__25823));
    InMux I__3175 (
            .O(N__25828),
            .I(N__25823));
    LocalMux I__3174 (
            .O(N__25823),
            .I(N__25820));
    Span12Mux_s10_v I__3173 (
            .O(N__25820),
            .I(N__25816));
    InMux I__3172 (
            .O(N__25819),
            .I(N__25813));
    Odrv12 I__3171 (
            .O(N__25816),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ));
    LocalMux I__3170 (
            .O(N__25813),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ));
    CascadeMux I__3169 (
            .O(N__25808),
            .I(N__25804));
    InMux I__3168 (
            .O(N__25807),
            .I(N__25801));
    InMux I__3167 (
            .O(N__25804),
            .I(N__25798));
    LocalMux I__3166 (
            .O(N__25801),
            .I(N__25795));
    LocalMux I__3165 (
            .O(N__25798),
            .I(N__25792));
    Span4Mux_v I__3164 (
            .O(N__25795),
            .I(N__25787));
    Span4Mux_v I__3163 (
            .O(N__25792),
            .I(N__25787));
    Odrv4 I__3162 (
            .O(N__25787),
            .I(\phase_controller_inst2.stoper_tr.counter ));
    InMux I__3161 (
            .O(N__25784),
            .I(N__25781));
    LocalMux I__3160 (
            .O(N__25781),
            .I(N__25778));
    Span4Mux_h I__3159 (
            .O(N__25778),
            .I(N__25775));
    Odrv4 I__3158 (
            .O(N__25775),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ));
    InMux I__3157 (
            .O(N__25772),
            .I(N__25768));
    InMux I__3156 (
            .O(N__25771),
            .I(N__25765));
    LocalMux I__3155 (
            .O(N__25768),
            .I(N__25762));
    LocalMux I__3154 (
            .O(N__25765),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ));
    Odrv12 I__3153 (
            .O(N__25762),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ));
    CascadeMux I__3152 (
            .O(N__25757),
            .I(N__25754));
    InMux I__3151 (
            .O(N__25754),
            .I(N__25751));
    LocalMux I__3150 (
            .O(N__25751),
            .I(\phase_controller_inst2.stoper_tr.counter_i_12 ));
    InMux I__3149 (
            .O(N__25748),
            .I(N__25744));
    InMux I__3148 (
            .O(N__25747),
            .I(N__25741));
    LocalMux I__3147 (
            .O(N__25744),
            .I(N__25738));
    LocalMux I__3146 (
            .O(N__25741),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ));
    Odrv12 I__3145 (
            .O(N__25738),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ));
    InMux I__3144 (
            .O(N__25733),
            .I(N__25730));
    LocalMux I__3143 (
            .O(N__25730),
            .I(N__25727));
    Span4Mux_v I__3142 (
            .O(N__25727),
            .I(N__25724));
    Odrv4 I__3141 (
            .O(N__25724),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ));
    CascadeMux I__3140 (
            .O(N__25721),
            .I(N__25718));
    InMux I__3139 (
            .O(N__25718),
            .I(N__25715));
    LocalMux I__3138 (
            .O(N__25715),
            .I(N__25712));
    Odrv4 I__3137 (
            .O(N__25712),
            .I(\phase_controller_inst2.stoper_tr.counter_i_13 ));
    InMux I__3136 (
            .O(N__25709),
            .I(N__25705));
    InMux I__3135 (
            .O(N__25708),
            .I(N__25702));
    LocalMux I__3134 (
            .O(N__25705),
            .I(N__25699));
    LocalMux I__3133 (
            .O(N__25702),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ));
    Odrv12 I__3132 (
            .O(N__25699),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ));
    InMux I__3131 (
            .O(N__25694),
            .I(N__25691));
    LocalMux I__3130 (
            .O(N__25691),
            .I(N__25688));
    Span4Mux_h I__3129 (
            .O(N__25688),
            .I(N__25685));
    Odrv4 I__3128 (
            .O(N__25685),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ));
    CascadeMux I__3127 (
            .O(N__25682),
            .I(N__25679));
    InMux I__3126 (
            .O(N__25679),
            .I(N__25676));
    LocalMux I__3125 (
            .O(N__25676),
            .I(\phase_controller_inst2.stoper_tr.counter_i_14 ));
    InMux I__3124 (
            .O(N__25673),
            .I(N__25670));
    LocalMux I__3123 (
            .O(N__25670),
            .I(N__25666));
    InMux I__3122 (
            .O(N__25669),
            .I(N__25663));
    Span4Mux_v I__3121 (
            .O(N__25666),
            .I(N__25660));
    LocalMux I__3120 (
            .O(N__25663),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ));
    Odrv4 I__3119 (
            .O(N__25660),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ));
    CascadeMux I__3118 (
            .O(N__25655),
            .I(N__25652));
    InMux I__3117 (
            .O(N__25652),
            .I(N__25649));
    LocalMux I__3116 (
            .O(N__25649),
            .I(N__25646));
    Span4Mux_v I__3115 (
            .O(N__25646),
            .I(N__25643));
    Odrv4 I__3114 (
            .O(N__25643),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ));
    InMux I__3113 (
            .O(N__25640),
            .I(N__25637));
    LocalMux I__3112 (
            .O(N__25637),
            .I(\phase_controller_inst2.stoper_tr.counter_i_15 ));
    InMux I__3111 (
            .O(N__25634),
            .I(N__25631));
    LocalMux I__3110 (
            .O(N__25631),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt16 ));
    CascadeMux I__3109 (
            .O(N__25628),
            .I(N__25625));
    InMux I__3108 (
            .O(N__25625),
            .I(N__25622));
    LocalMux I__3107 (
            .O(N__25622),
            .I(N__25619));
    Odrv4 I__3106 (
            .O(N__25619),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ));
    InMux I__3105 (
            .O(N__25616),
            .I(N__25613));
    LocalMux I__3104 (
            .O(N__25613),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ));
    CascadeMux I__3103 (
            .O(N__25610),
            .I(N__25607));
    InMux I__3102 (
            .O(N__25607),
            .I(N__25604));
    LocalMux I__3101 (
            .O(N__25604),
            .I(N__25601));
    Odrv4 I__3100 (
            .O(N__25601),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt18 ));
    InMux I__3099 (
            .O(N__25598),
            .I(N__25595));
    LocalMux I__3098 (
            .O(N__25595),
            .I(N__25592));
    Span4Mux_h I__3097 (
            .O(N__25592),
            .I(N__25589));
    Odrv4 I__3096 (
            .O(N__25589),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ));
    CascadeMux I__3095 (
            .O(N__25586),
            .I(N__25583));
    InMux I__3094 (
            .O(N__25583),
            .I(N__25580));
    LocalMux I__3093 (
            .O(N__25580),
            .I(N__25577));
    Span4Mux_v I__3092 (
            .O(N__25577),
            .I(N__25574));
    Odrv4 I__3091 (
            .O(N__25574),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt20 ));
    InMux I__3090 (
            .O(N__25571),
            .I(N__25568));
    LocalMux I__3089 (
            .O(N__25568),
            .I(N__25565));
    Odrv4 I__3088 (
            .O(N__25565),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ));
    CascadeMux I__3087 (
            .O(N__25562),
            .I(N__25559));
    InMux I__3086 (
            .O(N__25559),
            .I(N__25556));
    LocalMux I__3085 (
            .O(N__25556),
            .I(N__25553));
    Span4Mux_v I__3084 (
            .O(N__25553),
            .I(N__25550));
    Odrv4 I__3083 (
            .O(N__25550),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt22 ));
    InMux I__3082 (
            .O(N__25547),
            .I(N__25543));
    InMux I__3081 (
            .O(N__25546),
            .I(N__25540));
    LocalMux I__3080 (
            .O(N__25543),
            .I(N__25537));
    LocalMux I__3079 (
            .O(N__25540),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ));
    Odrv12 I__3078 (
            .O(N__25537),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ));
    InMux I__3077 (
            .O(N__25532),
            .I(N__25529));
    LocalMux I__3076 (
            .O(N__25529),
            .I(N__25526));
    Span4Mux_h I__3075 (
            .O(N__25526),
            .I(N__25523));
    Odrv4 I__3074 (
            .O(N__25523),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ));
    CascadeMux I__3073 (
            .O(N__25520),
            .I(N__25517));
    InMux I__3072 (
            .O(N__25517),
            .I(N__25514));
    LocalMux I__3071 (
            .O(N__25514),
            .I(\phase_controller_inst2.stoper_tr.counter_i_5 ));
    InMux I__3070 (
            .O(N__25511),
            .I(N__25508));
    LocalMux I__3069 (
            .O(N__25508),
            .I(N__25505));
    Span4Mux_v I__3068 (
            .O(N__25505),
            .I(N__25502));
    Odrv4 I__3067 (
            .O(N__25502),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ));
    InMux I__3066 (
            .O(N__25499),
            .I(N__25496));
    LocalMux I__3065 (
            .O(N__25496),
            .I(N__25492));
    InMux I__3064 (
            .O(N__25495),
            .I(N__25489));
    Span4Mux_v I__3063 (
            .O(N__25492),
            .I(N__25486));
    LocalMux I__3062 (
            .O(N__25489),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ));
    Odrv4 I__3061 (
            .O(N__25486),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ));
    CascadeMux I__3060 (
            .O(N__25481),
            .I(N__25478));
    InMux I__3059 (
            .O(N__25478),
            .I(N__25475));
    LocalMux I__3058 (
            .O(N__25475),
            .I(N__25472));
    Odrv4 I__3057 (
            .O(N__25472),
            .I(\phase_controller_inst2.stoper_tr.counter_i_6 ));
    InMux I__3056 (
            .O(N__25469),
            .I(N__25466));
    LocalMux I__3055 (
            .O(N__25466),
            .I(N__25463));
    Odrv4 I__3054 (
            .O(N__25463),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ));
    InMux I__3053 (
            .O(N__25460),
            .I(N__25457));
    LocalMux I__3052 (
            .O(N__25457),
            .I(N__25453));
    InMux I__3051 (
            .O(N__25456),
            .I(N__25450));
    Span4Mux_v I__3050 (
            .O(N__25453),
            .I(N__25447));
    LocalMux I__3049 (
            .O(N__25450),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ));
    Odrv4 I__3048 (
            .O(N__25447),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ));
    CascadeMux I__3047 (
            .O(N__25442),
            .I(N__25439));
    InMux I__3046 (
            .O(N__25439),
            .I(N__25436));
    LocalMux I__3045 (
            .O(N__25436),
            .I(\phase_controller_inst2.stoper_tr.counter_i_7 ));
    InMux I__3044 (
            .O(N__25433),
            .I(N__25429));
    InMux I__3043 (
            .O(N__25432),
            .I(N__25426));
    LocalMux I__3042 (
            .O(N__25429),
            .I(N__25423));
    LocalMux I__3041 (
            .O(N__25426),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ));
    Odrv12 I__3040 (
            .O(N__25423),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ));
    InMux I__3039 (
            .O(N__25418),
            .I(N__25415));
    LocalMux I__3038 (
            .O(N__25415),
            .I(N__25412));
    Span4Mux_v I__3037 (
            .O(N__25412),
            .I(N__25409));
    Odrv4 I__3036 (
            .O(N__25409),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ));
    CascadeMux I__3035 (
            .O(N__25406),
            .I(N__25403));
    InMux I__3034 (
            .O(N__25403),
            .I(N__25400));
    LocalMux I__3033 (
            .O(N__25400),
            .I(\phase_controller_inst2.stoper_tr.counter_i_8 ));
    InMux I__3032 (
            .O(N__25397),
            .I(N__25394));
    LocalMux I__3031 (
            .O(N__25394),
            .I(N__25391));
    Span4Mux_v I__3030 (
            .O(N__25391),
            .I(N__25388));
    Odrv4 I__3029 (
            .O(N__25388),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ));
    InMux I__3028 (
            .O(N__25385),
            .I(N__25381));
    InMux I__3027 (
            .O(N__25384),
            .I(N__25378));
    LocalMux I__3026 (
            .O(N__25381),
            .I(N__25375));
    LocalMux I__3025 (
            .O(N__25378),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ));
    Odrv12 I__3024 (
            .O(N__25375),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ));
    CascadeMux I__3023 (
            .O(N__25370),
            .I(N__25367));
    InMux I__3022 (
            .O(N__25367),
            .I(N__25364));
    LocalMux I__3021 (
            .O(N__25364),
            .I(\phase_controller_inst2.stoper_tr.counter_i_9 ));
    InMux I__3020 (
            .O(N__25361),
            .I(N__25358));
    LocalMux I__3019 (
            .O(N__25358),
            .I(N__25355));
    Span4Mux_h I__3018 (
            .O(N__25355),
            .I(N__25352));
    Odrv4 I__3017 (
            .O(N__25352),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ));
    InMux I__3016 (
            .O(N__25349),
            .I(N__25345));
    InMux I__3015 (
            .O(N__25348),
            .I(N__25342));
    LocalMux I__3014 (
            .O(N__25345),
            .I(N__25339));
    LocalMux I__3013 (
            .O(N__25342),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ));
    Odrv12 I__3012 (
            .O(N__25339),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ));
    CascadeMux I__3011 (
            .O(N__25334),
            .I(N__25331));
    InMux I__3010 (
            .O(N__25331),
            .I(N__25328));
    LocalMux I__3009 (
            .O(N__25328),
            .I(\phase_controller_inst2.stoper_tr.counter_i_10 ));
    CascadeMux I__3008 (
            .O(N__25325),
            .I(N__25322));
    InMux I__3007 (
            .O(N__25322),
            .I(N__25319));
    LocalMux I__3006 (
            .O(N__25319),
            .I(N__25316));
    Odrv4 I__3005 (
            .O(N__25316),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ));
    InMux I__3004 (
            .O(N__25313),
            .I(N__25309));
    InMux I__3003 (
            .O(N__25312),
            .I(N__25306));
    LocalMux I__3002 (
            .O(N__25309),
            .I(N__25303));
    LocalMux I__3001 (
            .O(N__25306),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ));
    Odrv12 I__3000 (
            .O(N__25303),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ));
    InMux I__2999 (
            .O(N__25298),
            .I(N__25295));
    LocalMux I__2998 (
            .O(N__25295),
            .I(\phase_controller_inst2.stoper_tr.counter_i_11 ));
    InMux I__2997 (
            .O(N__25292),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_28 ));
    InMux I__2996 (
            .O(N__25289),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_29 ));
    InMux I__2995 (
            .O(N__25286),
            .I(N__25246));
    InMux I__2994 (
            .O(N__25285),
            .I(N__25246));
    InMux I__2993 (
            .O(N__25284),
            .I(N__25246));
    InMux I__2992 (
            .O(N__25283),
            .I(N__25246));
    InMux I__2991 (
            .O(N__25282),
            .I(N__25237));
    InMux I__2990 (
            .O(N__25281),
            .I(N__25237));
    InMux I__2989 (
            .O(N__25280),
            .I(N__25237));
    InMux I__2988 (
            .O(N__25279),
            .I(N__25237));
    InMux I__2987 (
            .O(N__25278),
            .I(N__25228));
    InMux I__2986 (
            .O(N__25277),
            .I(N__25228));
    InMux I__2985 (
            .O(N__25276),
            .I(N__25228));
    InMux I__2984 (
            .O(N__25275),
            .I(N__25228));
    InMux I__2983 (
            .O(N__25274),
            .I(N__25219));
    InMux I__2982 (
            .O(N__25273),
            .I(N__25219));
    InMux I__2981 (
            .O(N__25272),
            .I(N__25219));
    InMux I__2980 (
            .O(N__25271),
            .I(N__25219));
    InMux I__2979 (
            .O(N__25270),
            .I(N__25210));
    InMux I__2978 (
            .O(N__25269),
            .I(N__25210));
    InMux I__2977 (
            .O(N__25268),
            .I(N__25210));
    InMux I__2976 (
            .O(N__25267),
            .I(N__25210));
    InMux I__2975 (
            .O(N__25266),
            .I(N__25201));
    InMux I__2974 (
            .O(N__25265),
            .I(N__25201));
    InMux I__2973 (
            .O(N__25264),
            .I(N__25201));
    InMux I__2972 (
            .O(N__25263),
            .I(N__25201));
    InMux I__2971 (
            .O(N__25262),
            .I(N__25192));
    InMux I__2970 (
            .O(N__25261),
            .I(N__25192));
    InMux I__2969 (
            .O(N__25260),
            .I(N__25192));
    InMux I__2968 (
            .O(N__25259),
            .I(N__25192));
    InMux I__2967 (
            .O(N__25258),
            .I(N__25183));
    InMux I__2966 (
            .O(N__25257),
            .I(N__25183));
    InMux I__2965 (
            .O(N__25256),
            .I(N__25183));
    InMux I__2964 (
            .O(N__25255),
            .I(N__25183));
    LocalMux I__2963 (
            .O(N__25246),
            .I(N__25176));
    LocalMux I__2962 (
            .O(N__25237),
            .I(N__25176));
    LocalMux I__2961 (
            .O(N__25228),
            .I(N__25176));
    LocalMux I__2960 (
            .O(N__25219),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    LocalMux I__2959 (
            .O(N__25210),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    LocalMux I__2958 (
            .O(N__25201),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    LocalMux I__2957 (
            .O(N__25192),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    LocalMux I__2956 (
            .O(N__25183),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    Odrv4 I__2955 (
            .O(N__25176),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    InMux I__2954 (
            .O(N__25163),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_30 ));
    CEMux I__2953 (
            .O(N__25160),
            .I(N__25148));
    CEMux I__2952 (
            .O(N__25159),
            .I(N__25148));
    CEMux I__2951 (
            .O(N__25158),
            .I(N__25148));
    CEMux I__2950 (
            .O(N__25157),
            .I(N__25148));
    GlobalMux I__2949 (
            .O(N__25148),
            .I(N__25145));
    gio2CtrlBuf I__2948 (
            .O(N__25145),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0_g ));
    InMux I__2947 (
            .O(N__25142),
            .I(N__25139));
    LocalMux I__2946 (
            .O(N__25139),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ));
    InMux I__2945 (
            .O(N__25136),
            .I(N__25132));
    InMux I__2944 (
            .O(N__25135),
            .I(N__25129));
    LocalMux I__2943 (
            .O(N__25132),
            .I(N__25126));
    LocalMux I__2942 (
            .O(N__25129),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ));
    Odrv12 I__2941 (
            .O(N__25126),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ));
    CascadeMux I__2940 (
            .O(N__25121),
            .I(N__25118));
    InMux I__2939 (
            .O(N__25118),
            .I(N__25115));
    LocalMux I__2938 (
            .O(N__25115),
            .I(\phase_controller_inst2.stoper_tr.counter_i_0 ));
    InMux I__2937 (
            .O(N__25112),
            .I(N__25109));
    LocalMux I__2936 (
            .O(N__25109),
            .I(N__25106));
    Odrv4 I__2935 (
            .O(N__25106),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ));
    InMux I__2934 (
            .O(N__25103),
            .I(N__25099));
    InMux I__2933 (
            .O(N__25102),
            .I(N__25096));
    LocalMux I__2932 (
            .O(N__25099),
            .I(N__25093));
    LocalMux I__2931 (
            .O(N__25096),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ));
    Odrv12 I__2930 (
            .O(N__25093),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ));
    CascadeMux I__2929 (
            .O(N__25088),
            .I(N__25085));
    InMux I__2928 (
            .O(N__25085),
            .I(N__25082));
    LocalMux I__2927 (
            .O(N__25082),
            .I(\phase_controller_inst2.stoper_tr.counter_i_1 ));
    InMux I__2926 (
            .O(N__25079),
            .I(N__25076));
    LocalMux I__2925 (
            .O(N__25076),
            .I(N__25073));
    Span4Mux_h I__2924 (
            .O(N__25073),
            .I(N__25070));
    Odrv4 I__2923 (
            .O(N__25070),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ));
    InMux I__2922 (
            .O(N__25067),
            .I(N__25063));
    InMux I__2921 (
            .O(N__25066),
            .I(N__25060));
    LocalMux I__2920 (
            .O(N__25063),
            .I(N__25057));
    LocalMux I__2919 (
            .O(N__25060),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ));
    Odrv12 I__2918 (
            .O(N__25057),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ));
    CascadeMux I__2917 (
            .O(N__25052),
            .I(N__25049));
    InMux I__2916 (
            .O(N__25049),
            .I(N__25046));
    LocalMux I__2915 (
            .O(N__25046),
            .I(N__25043));
    Odrv4 I__2914 (
            .O(N__25043),
            .I(\phase_controller_inst2.stoper_tr.counter_i_2 ));
    InMux I__2913 (
            .O(N__25040),
            .I(N__25037));
    LocalMux I__2912 (
            .O(N__25037),
            .I(N__25034));
    Span4Mux_h I__2911 (
            .O(N__25034),
            .I(N__25031));
    Odrv4 I__2910 (
            .O(N__25031),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ));
    InMux I__2909 (
            .O(N__25028),
            .I(N__25024));
    InMux I__2908 (
            .O(N__25027),
            .I(N__25021));
    LocalMux I__2907 (
            .O(N__25024),
            .I(N__25018));
    LocalMux I__2906 (
            .O(N__25021),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ));
    Odrv12 I__2905 (
            .O(N__25018),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ));
    CascadeMux I__2904 (
            .O(N__25013),
            .I(N__25010));
    InMux I__2903 (
            .O(N__25010),
            .I(N__25007));
    LocalMux I__2902 (
            .O(N__25007),
            .I(\phase_controller_inst2.stoper_tr.counter_i_3 ));
    InMux I__2901 (
            .O(N__25004),
            .I(N__25001));
    LocalMux I__2900 (
            .O(N__25001),
            .I(N__24998));
    Span4Mux_h I__2899 (
            .O(N__24998),
            .I(N__24995));
    Odrv4 I__2898 (
            .O(N__24995),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ));
    InMux I__2897 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__2896 (
            .O(N__24989),
            .I(N__24985));
    InMux I__2895 (
            .O(N__24988),
            .I(N__24982));
    Span4Mux_v I__2894 (
            .O(N__24985),
            .I(N__24979));
    LocalMux I__2893 (
            .O(N__24982),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ));
    Odrv4 I__2892 (
            .O(N__24979),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ));
    CascadeMux I__2891 (
            .O(N__24974),
            .I(N__24971));
    InMux I__2890 (
            .O(N__24971),
            .I(N__24968));
    LocalMux I__2889 (
            .O(N__24968),
            .I(N__24965));
    Odrv4 I__2888 (
            .O(N__24965),
            .I(\phase_controller_inst2.stoper_tr.counter_i_4 ));
    InMux I__2887 (
            .O(N__24962),
            .I(N__24957));
    InMux I__2886 (
            .O(N__24961),
            .I(N__24952));
    InMux I__2885 (
            .O(N__24960),
            .I(N__24952));
    LocalMux I__2884 (
            .O(N__24957),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ));
    LocalMux I__2883 (
            .O(N__24952),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ));
    InMux I__2882 (
            .O(N__24947),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_20 ));
    InMux I__2881 (
            .O(N__24944),
            .I(N__24939));
    InMux I__2880 (
            .O(N__24943),
            .I(N__24934));
    InMux I__2879 (
            .O(N__24942),
            .I(N__24934));
    LocalMux I__2878 (
            .O(N__24939),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_22 ));
    LocalMux I__2877 (
            .O(N__24934),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_22 ));
    InMux I__2876 (
            .O(N__24929),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_21 ));
    InMux I__2875 (
            .O(N__24926),
            .I(N__24921));
    InMux I__2874 (
            .O(N__24925),
            .I(N__24916));
    InMux I__2873 (
            .O(N__24924),
            .I(N__24916));
    LocalMux I__2872 (
            .O(N__24921),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_23 ));
    LocalMux I__2871 (
            .O(N__24916),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_23 ));
    InMux I__2870 (
            .O(N__24911),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_22 ));
    InMux I__2869 (
            .O(N__24908),
            .I(N__24903));
    InMux I__2868 (
            .O(N__24907),
            .I(N__24898));
    InMux I__2867 (
            .O(N__24906),
            .I(N__24898));
    LocalMux I__2866 (
            .O(N__24903),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ));
    LocalMux I__2865 (
            .O(N__24898),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ));
    InMux I__2864 (
            .O(N__24893),
            .I(bfn_8_11_0_));
    InMux I__2863 (
            .O(N__24890),
            .I(N__24885));
    InMux I__2862 (
            .O(N__24889),
            .I(N__24880));
    InMux I__2861 (
            .O(N__24888),
            .I(N__24880));
    LocalMux I__2860 (
            .O(N__24885),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ));
    LocalMux I__2859 (
            .O(N__24880),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ));
    InMux I__2858 (
            .O(N__24875),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_24 ));
    InMux I__2857 (
            .O(N__24872),
            .I(N__24867));
    InMux I__2856 (
            .O(N__24871),
            .I(N__24862));
    InMux I__2855 (
            .O(N__24870),
            .I(N__24862));
    LocalMux I__2854 (
            .O(N__24867),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ));
    LocalMux I__2853 (
            .O(N__24862),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ));
    InMux I__2852 (
            .O(N__24857),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_25 ));
    CascadeMux I__2851 (
            .O(N__24854),
            .I(N__24849));
    CascadeMux I__2850 (
            .O(N__24853),
            .I(N__24846));
    InMux I__2849 (
            .O(N__24852),
            .I(N__24843));
    InMux I__2848 (
            .O(N__24849),
            .I(N__24838));
    InMux I__2847 (
            .O(N__24846),
            .I(N__24838));
    LocalMux I__2846 (
            .O(N__24843),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ));
    LocalMux I__2845 (
            .O(N__24838),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ));
    InMux I__2844 (
            .O(N__24833),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_26 ));
    InMux I__2843 (
            .O(N__24830),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_27 ));
    InMux I__2842 (
            .O(N__24827),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_11 ));
    InMux I__2841 (
            .O(N__24824),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_12 ));
    InMux I__2840 (
            .O(N__24821),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_13 ));
    InMux I__2839 (
            .O(N__24818),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_14 ));
    CascadeMux I__2838 (
            .O(N__24815),
            .I(N__24811));
    CascadeMux I__2837 (
            .O(N__24814),
            .I(N__24808));
    InMux I__2836 (
            .O(N__24811),
            .I(N__24803));
    InMux I__2835 (
            .O(N__24808),
            .I(N__24803));
    LocalMux I__2834 (
            .O(N__24803),
            .I(N__24799));
    InMux I__2833 (
            .O(N__24802),
            .I(N__24796));
    Span4Mux_v I__2832 (
            .O(N__24799),
            .I(N__24793));
    LocalMux I__2831 (
            .O(N__24796),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ));
    Odrv4 I__2830 (
            .O(N__24793),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ));
    InMux I__2829 (
            .O(N__24788),
            .I(bfn_8_10_0_));
    InMux I__2828 (
            .O(N__24785),
            .I(N__24779));
    InMux I__2827 (
            .O(N__24784),
            .I(N__24779));
    LocalMux I__2826 (
            .O(N__24779),
            .I(N__24775));
    InMux I__2825 (
            .O(N__24778),
            .I(N__24772));
    Span4Mux_v I__2824 (
            .O(N__24775),
            .I(N__24769));
    LocalMux I__2823 (
            .O(N__24772),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ));
    Odrv4 I__2822 (
            .O(N__24769),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ));
    InMux I__2821 (
            .O(N__24764),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_16 ));
    CascadeMux I__2820 (
            .O(N__24761),
            .I(N__24757));
    CascadeMux I__2819 (
            .O(N__24760),
            .I(N__24754));
    InMux I__2818 (
            .O(N__24757),
            .I(N__24749));
    InMux I__2817 (
            .O(N__24754),
            .I(N__24749));
    LocalMux I__2816 (
            .O(N__24749),
            .I(N__24745));
    InMux I__2815 (
            .O(N__24748),
            .I(N__24742));
    Span4Mux_v I__2814 (
            .O(N__24745),
            .I(N__24739));
    LocalMux I__2813 (
            .O(N__24742),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ));
    Odrv4 I__2812 (
            .O(N__24739),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ));
    InMux I__2811 (
            .O(N__24734),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_17 ));
    InMux I__2810 (
            .O(N__24731),
            .I(N__24725));
    InMux I__2809 (
            .O(N__24730),
            .I(N__24725));
    LocalMux I__2808 (
            .O(N__24725),
            .I(N__24721));
    InMux I__2807 (
            .O(N__24724),
            .I(N__24718));
    Span4Mux_v I__2806 (
            .O(N__24721),
            .I(N__24715));
    LocalMux I__2805 (
            .O(N__24718),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ));
    Odrv4 I__2804 (
            .O(N__24715),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ));
    InMux I__2803 (
            .O(N__24710),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_18 ));
    InMux I__2802 (
            .O(N__24707),
            .I(N__24702));
    InMux I__2801 (
            .O(N__24706),
            .I(N__24697));
    InMux I__2800 (
            .O(N__24705),
            .I(N__24697));
    LocalMux I__2799 (
            .O(N__24702),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ));
    LocalMux I__2798 (
            .O(N__24697),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ));
    InMux I__2797 (
            .O(N__24692),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_19 ));
    InMux I__2796 (
            .O(N__24689),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_2 ));
    InMux I__2795 (
            .O(N__24686),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_3 ));
    InMux I__2794 (
            .O(N__24683),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_4 ));
    InMux I__2793 (
            .O(N__24680),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_5 ));
    InMux I__2792 (
            .O(N__24677),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_6 ));
    InMux I__2791 (
            .O(N__24674),
            .I(bfn_8_9_0_));
    InMux I__2790 (
            .O(N__24671),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_8 ));
    InMux I__2789 (
            .O(N__24668),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_9 ));
    InMux I__2788 (
            .O(N__24665),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_10 ));
    CascadeMux I__2787 (
            .O(N__24662),
            .I(N__24659));
    InMux I__2786 (
            .O(N__24659),
            .I(N__24656));
    LocalMux I__2785 (
            .O(N__24656),
            .I(\phase_controller_inst2.stoper_tr.un4_start_0 ));
    InMux I__2784 (
            .O(N__24653),
            .I(N__24644));
    InMux I__2783 (
            .O(N__24652),
            .I(N__24644));
    InMux I__2782 (
            .O(N__24651),
            .I(N__24644));
    LocalMux I__2781 (
            .O(N__24644),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    CascadeMux I__2780 (
            .O(N__24641),
            .I(N__24636));
    CascadeMux I__2779 (
            .O(N__24640),
            .I(N__24633));
    InMux I__2778 (
            .O(N__24639),
            .I(N__24626));
    InMux I__2777 (
            .O(N__24636),
            .I(N__24626));
    InMux I__2776 (
            .O(N__24633),
            .I(N__24626));
    LocalMux I__2775 (
            .O(N__24626),
            .I(\phase_controller_inst2.start_flagZ0 ));
    InMux I__2774 (
            .O(N__24623),
            .I(N__24616));
    InMux I__2773 (
            .O(N__24622),
            .I(N__24612));
    InMux I__2772 (
            .O(N__24621),
            .I(N__24607));
    InMux I__2771 (
            .O(N__24620),
            .I(N__24607));
    InMux I__2770 (
            .O(N__24619),
            .I(N__24604));
    LocalMux I__2769 (
            .O(N__24616),
            .I(N__24601));
    InMux I__2768 (
            .O(N__24615),
            .I(N__24598));
    LocalMux I__2767 (
            .O(N__24612),
            .I(N__24595));
    LocalMux I__2766 (
            .O(N__24607),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__2765 (
            .O(N__24604),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__2764 (
            .O(N__24601),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__2763 (
            .O(N__24598),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__2762 (
            .O(N__24595),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__2761 (
            .O(N__24584),
            .I(N__24577));
    InMux I__2760 (
            .O(N__24583),
            .I(N__24577));
    InMux I__2759 (
            .O(N__24582),
            .I(N__24574));
    LocalMux I__2758 (
            .O(N__24577),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    LocalMux I__2757 (
            .O(N__24574),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__2756 (
            .O(N__24569),
            .I(N__24566));
    LocalMux I__2755 (
            .O(N__24566),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    InMux I__2754 (
            .O(N__24563),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_0 ));
    InMux I__2753 (
            .O(N__24560),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_1 ));
    InMux I__2752 (
            .O(N__24557),
            .I(N__24551));
    InMux I__2751 (
            .O(N__24556),
            .I(N__24551));
    LocalMux I__2750 (
            .O(N__24551),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ));
    InMux I__2749 (
            .O(N__24548),
            .I(N__24542));
    InMux I__2748 (
            .O(N__24547),
            .I(N__24542));
    LocalMux I__2747 (
            .O(N__24542),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ));
    IoInMux I__2746 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__2745 (
            .O(N__24536),
            .I(N__24533));
    Span4Mux_s1_v I__2744 (
            .O(N__24533),
            .I(N__24530));
    Span4Mux_h I__2743 (
            .O(N__24530),
            .I(N__24527));
    Odrv4 I__2742 (
            .O(N__24527),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__2741 (
            .O(N__24524),
            .I(N__24518));
    InMux I__2740 (
            .O(N__24523),
            .I(N__24518));
    LocalMux I__2739 (
            .O(N__24518),
            .I(N__24515));
    Odrv12 I__2738 (
            .O(N__24515),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ));
    InMux I__2737 (
            .O(N__24512),
            .I(N__24506));
    InMux I__2736 (
            .O(N__24511),
            .I(N__24506));
    LocalMux I__2735 (
            .O(N__24506),
            .I(N__24503));
    Span12Mux_v I__2734 (
            .O(N__24503),
            .I(N__24500));
    Odrv12 I__2733 (
            .O(N__24500),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ));
    InMux I__2732 (
            .O(N__24497),
            .I(N__24491));
    InMux I__2731 (
            .O(N__24496),
            .I(N__24491));
    LocalMux I__2730 (
            .O(N__24491),
            .I(N__24488));
    Odrv12 I__2729 (
            .O(N__24488),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ));
    CascadeMux I__2728 (
            .O(N__24485),
            .I(N__24481));
    CascadeMux I__2727 (
            .O(N__24484),
            .I(N__24478));
    InMux I__2726 (
            .O(N__24481),
            .I(N__24473));
    InMux I__2725 (
            .O(N__24478),
            .I(N__24473));
    LocalMux I__2724 (
            .O(N__24473),
            .I(N__24470));
    Span4Mux_v I__2723 (
            .O(N__24470),
            .I(N__24467));
    Span4Mux_v I__2722 (
            .O(N__24467),
            .I(N__24464));
    Odrv4 I__2721 (
            .O(N__24464),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ));
    CEMux I__2720 (
            .O(N__24461),
            .I(N__24458));
    LocalMux I__2719 (
            .O(N__24458),
            .I(N__24452));
    CEMux I__2718 (
            .O(N__24457),
            .I(N__24449));
    CEMux I__2717 (
            .O(N__24456),
            .I(N__24444));
    CEMux I__2716 (
            .O(N__24455),
            .I(N__24440));
    Span4Mux_v I__2715 (
            .O(N__24452),
            .I(N__24432));
    LocalMux I__2714 (
            .O(N__24449),
            .I(N__24432));
    CEMux I__2713 (
            .O(N__24448),
            .I(N__24429));
    CEMux I__2712 (
            .O(N__24447),
            .I(N__24426));
    LocalMux I__2711 (
            .O(N__24444),
            .I(N__24423));
    CEMux I__2710 (
            .O(N__24443),
            .I(N__24420));
    LocalMux I__2709 (
            .O(N__24440),
            .I(N__24417));
    CEMux I__2708 (
            .O(N__24439),
            .I(N__24414));
    CEMux I__2707 (
            .O(N__24438),
            .I(N__24411));
    CEMux I__2706 (
            .O(N__24437),
            .I(N__24408));
    Span4Mux_h I__2705 (
            .O(N__24432),
            .I(N__24401));
    LocalMux I__2704 (
            .O(N__24429),
            .I(N__24401));
    LocalMux I__2703 (
            .O(N__24426),
            .I(N__24398));
    Span4Mux_h I__2702 (
            .O(N__24423),
            .I(N__24395));
    LocalMux I__2701 (
            .O(N__24420),
            .I(N__24392));
    Span4Mux_h I__2700 (
            .O(N__24417),
            .I(N__24387));
    LocalMux I__2699 (
            .O(N__24414),
            .I(N__24387));
    LocalMux I__2698 (
            .O(N__24411),
            .I(N__24382));
    LocalMux I__2697 (
            .O(N__24408),
            .I(N__24382));
    CEMux I__2696 (
            .O(N__24407),
            .I(N__24379));
    CEMux I__2695 (
            .O(N__24406),
            .I(N__24376));
    Span4Mux_v I__2694 (
            .O(N__24401),
            .I(N__24373));
    Span4Mux_v I__2693 (
            .O(N__24398),
            .I(N__24370));
    Span4Mux_h I__2692 (
            .O(N__24395),
            .I(N__24365));
    Span4Mux_h I__2691 (
            .O(N__24392),
            .I(N__24365));
    Span4Mux_v I__2690 (
            .O(N__24387),
            .I(N__24356));
    Span4Mux_v I__2689 (
            .O(N__24382),
            .I(N__24356));
    LocalMux I__2688 (
            .O(N__24379),
            .I(N__24356));
    LocalMux I__2687 (
            .O(N__24376),
            .I(N__24356));
    Span4Mux_h I__2686 (
            .O(N__24373),
            .I(N__24353));
    Span4Mux_v I__2685 (
            .O(N__24370),
            .I(N__24350));
    Span4Mux_v I__2684 (
            .O(N__24365),
            .I(N__24347));
    Span4Mux_v I__2683 (
            .O(N__24356),
            .I(N__24344));
    Odrv4 I__2682 (
            .O(N__24353),
            .I(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv4 I__2681 (
            .O(N__24350),
            .I(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv4 I__2680 (
            .O(N__24347),
            .I(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv4 I__2679 (
            .O(N__24344),
            .I(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ));
    InMux I__2678 (
            .O(N__24335),
            .I(N__24329));
    InMux I__2677 (
            .O(N__24334),
            .I(N__24329));
    LocalMux I__2676 (
            .O(N__24329),
            .I(N__24326));
    Odrv12 I__2675 (
            .O(N__24326),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ));
    CascadeMux I__2674 (
            .O(N__24323),
            .I(N__24319));
    CascadeMux I__2673 (
            .O(N__24322),
            .I(N__24316));
    InMux I__2672 (
            .O(N__24319),
            .I(N__24311));
    InMux I__2671 (
            .O(N__24316),
            .I(N__24311));
    LocalMux I__2670 (
            .O(N__24311),
            .I(N__24308));
    Odrv12 I__2669 (
            .O(N__24308),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ));
    InMux I__2668 (
            .O(N__24305),
            .I(N__24299));
    InMux I__2667 (
            .O(N__24304),
            .I(N__24299));
    LocalMux I__2666 (
            .O(N__24299),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ));
    InMux I__2665 (
            .O(N__24296),
            .I(N__24290));
    InMux I__2664 (
            .O(N__24295),
            .I(N__24290));
    LocalMux I__2663 (
            .O(N__24290),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ));
    InMux I__2662 (
            .O(N__24287),
            .I(N__24281));
    InMux I__2661 (
            .O(N__24286),
            .I(N__24281));
    LocalMux I__2660 (
            .O(N__24281),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ));
    InMux I__2659 (
            .O(N__24278),
            .I(N__24272));
    InMux I__2658 (
            .O(N__24277),
            .I(N__24272));
    LocalMux I__2657 (
            .O(N__24272),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ));
    CascadeMux I__2656 (
            .O(N__24269),
            .I(N__24265));
    CascadeMux I__2655 (
            .O(N__24268),
            .I(N__24262));
    InMux I__2654 (
            .O(N__24265),
            .I(N__24257));
    InMux I__2653 (
            .O(N__24262),
            .I(N__24257));
    LocalMux I__2652 (
            .O(N__24257),
            .I(N__24254));
    Span4Mux_h I__2651 (
            .O(N__24254),
            .I(N__24251));
    Span4Mux_v I__2650 (
            .O(N__24251),
            .I(N__24248));
    Odrv4 I__2649 (
            .O(N__24248),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ));
    CascadeMux I__2648 (
            .O(N__24245),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31_cascade_));
    InMux I__2647 (
            .O(N__24242),
            .I(N__24239));
    LocalMux I__2646 (
            .O(N__24239),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    CascadeMux I__2645 (
            .O(N__24236),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_));
    InMux I__2644 (
            .O(N__24233),
            .I(N__24227));
    InMux I__2643 (
            .O(N__24232),
            .I(N__24227));
    LocalMux I__2642 (
            .O(N__24227),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ));
    InMux I__2641 (
            .O(N__24224),
            .I(N__24219));
    InMux I__2640 (
            .O(N__24223),
            .I(N__24216));
    InMux I__2639 (
            .O(N__24222),
            .I(N__24213));
    LocalMux I__2638 (
            .O(N__24219),
            .I(N__24210));
    LocalMux I__2637 (
            .O(N__24216),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2636 (
            .O(N__24213),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__2635 (
            .O(N__24210),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    CascadeMux I__2634 (
            .O(N__24203),
            .I(N__24200));
    InMux I__2633 (
            .O(N__24200),
            .I(N__24197));
    LocalMux I__2632 (
            .O(N__24197),
            .I(N__24194));
    Odrv4 I__2631 (
            .O(N__24194),
            .I(\pwm_generator_inst.N_184_i ));
    InMux I__2630 (
            .O(N__24191),
            .I(N__24188));
    LocalMux I__2629 (
            .O(N__24188),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__2628 (
            .O(N__24185),
            .I(N__24180));
    InMux I__2627 (
            .O(N__24184),
            .I(N__24177));
    InMux I__2626 (
            .O(N__24183),
            .I(N__24174));
    LocalMux I__2625 (
            .O(N__24180),
            .I(N__24171));
    LocalMux I__2624 (
            .O(N__24177),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2623 (
            .O(N__24174),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__2622 (
            .O(N__24171),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    CascadeMux I__2621 (
            .O(N__24164),
            .I(N__24161));
    InMux I__2620 (
            .O(N__24161),
            .I(N__24158));
    LocalMux I__2619 (
            .O(N__24158),
            .I(N__24155));
    Span4Mux_h I__2618 (
            .O(N__24155),
            .I(N__24152));
    Odrv4 I__2617 (
            .O(N__24152),
            .I(\pwm_generator_inst.N_185_i ));
    InMux I__2616 (
            .O(N__24149),
            .I(N__24146));
    LocalMux I__2615 (
            .O(N__24146),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2614 (
            .O(N__24143),
            .I(N__24140));
    InMux I__2613 (
            .O(N__24140),
            .I(N__24137));
    LocalMux I__2612 (
            .O(N__24137),
            .I(N__24134));
    Span4Mux_v I__2611 (
            .O(N__24134),
            .I(N__24131));
    Odrv4 I__2610 (
            .O(N__24131),
            .I(\pwm_generator_inst.N_186_i ));
    InMux I__2609 (
            .O(N__24128),
            .I(N__24123));
    InMux I__2608 (
            .O(N__24127),
            .I(N__24120));
    InMux I__2607 (
            .O(N__24126),
            .I(N__24117));
    LocalMux I__2606 (
            .O(N__24123),
            .I(N__24114));
    LocalMux I__2605 (
            .O(N__24120),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2604 (
            .O(N__24117),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2603 (
            .O(N__24114),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2602 (
            .O(N__24107),
            .I(N__24104));
    LocalMux I__2601 (
            .O(N__24104),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2600 (
            .O(N__24101),
            .I(N__24098));
    InMux I__2599 (
            .O(N__24098),
            .I(N__24095));
    LocalMux I__2598 (
            .O(N__24095),
            .I(\pwm_generator_inst.N_187_i ));
    InMux I__2597 (
            .O(N__24092),
            .I(N__24088));
    InMux I__2596 (
            .O(N__24091),
            .I(N__24084));
    LocalMux I__2595 (
            .O(N__24088),
            .I(N__24081));
    InMux I__2594 (
            .O(N__24087),
            .I(N__24078));
    LocalMux I__2593 (
            .O(N__24084),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv12 I__2592 (
            .O(N__24081),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2591 (
            .O(N__24078),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2590 (
            .O(N__24071),
            .I(N__24068));
    LocalMux I__2589 (
            .O(N__24068),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__2588 (
            .O(N__24065),
            .I(N__24062));
    InMux I__2587 (
            .O(N__24062),
            .I(N__24059));
    LocalMux I__2586 (
            .O(N__24059),
            .I(N__24056));
    Odrv4 I__2585 (
            .O(N__24056),
            .I(\pwm_generator_inst.N_188_i ));
    InMux I__2584 (
            .O(N__24053),
            .I(N__24049));
    InMux I__2583 (
            .O(N__24052),
            .I(N__24045));
    LocalMux I__2582 (
            .O(N__24049),
            .I(N__24042));
    InMux I__2581 (
            .O(N__24048),
            .I(N__24039));
    LocalMux I__2580 (
            .O(N__24045),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv12 I__2579 (
            .O(N__24042),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2578 (
            .O(N__24039),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__2577 (
            .O(N__24032),
            .I(N__24029));
    LocalMux I__2576 (
            .O(N__24029),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2575 (
            .O(N__24026),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2574 (
            .O(N__24023),
            .I(N__24020));
    LocalMux I__2573 (
            .O(N__24020),
            .I(N__24017));
    Span4Mux_s3_v I__2572 (
            .O(N__24017),
            .I(N__24014));
    Sp12to4 I__2571 (
            .O(N__24014),
            .I(N__24011));
    Span12Mux_h I__2570 (
            .O(N__24011),
            .I(N__24008));
    Span12Mux_v I__2569 (
            .O(N__24008),
            .I(N__24005));
    Odrv12 I__2568 (
            .O(N__24005),
            .I(pwm_output_c));
    InMux I__2567 (
            .O(N__24002),
            .I(N__23999));
    LocalMux I__2566 (
            .O(N__23999),
            .I(N__23995));
    CascadeMux I__2565 (
            .O(N__23998),
            .I(N__23992));
    Span4Mux_h I__2564 (
            .O(N__23995),
            .I(N__23989));
    InMux I__2563 (
            .O(N__23992),
            .I(N__23986));
    Odrv4 I__2562 (
            .O(N__23989),
            .I(\pwm_generator_inst.un18_threshold1_20 ));
    LocalMux I__2561 (
            .O(N__23986),
            .I(\pwm_generator_inst.un18_threshold1_20 ));
    InMux I__2560 (
            .O(N__23981),
            .I(N__23978));
    LocalMux I__2559 (
            .O(N__23978),
            .I(\pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO ));
    CascadeMux I__2558 (
            .O(N__23975),
            .I(N__23972));
    InMux I__2557 (
            .O(N__23972),
            .I(N__23969));
    LocalMux I__2556 (
            .O(N__23969),
            .I(N__23966));
    Span4Mux_v I__2555 (
            .O(N__23966),
            .I(N__23962));
    InMux I__2554 (
            .O(N__23965),
            .I(N__23959));
    Odrv4 I__2553 (
            .O(N__23962),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0 ));
    LocalMux I__2552 (
            .O(N__23959),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0 ));
    InMux I__2551 (
            .O(N__23954),
            .I(N__23951));
    LocalMux I__2550 (
            .O(N__23951),
            .I(\pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO ));
    CascadeMux I__2549 (
            .O(N__23948),
            .I(N__23945));
    InMux I__2548 (
            .O(N__23945),
            .I(N__23942));
    LocalMux I__2547 (
            .O(N__23942),
            .I(N__23939));
    Span4Mux_h I__2546 (
            .O(N__23939),
            .I(N__23935));
    InMux I__2545 (
            .O(N__23938),
            .I(N__23932));
    Odrv4 I__2544 (
            .O(N__23935),
            .I(\pwm_generator_inst.un18_threshold1_21 ));
    LocalMux I__2543 (
            .O(N__23932),
            .I(\pwm_generator_inst.un18_threshold1_21 ));
    InMux I__2542 (
            .O(N__23927),
            .I(N__23924));
    LocalMux I__2541 (
            .O(N__23924),
            .I(N__23921));
    Span4Mux_h I__2540 (
            .O(N__23921),
            .I(N__23917));
    InMux I__2539 (
            .O(N__23920),
            .I(N__23914));
    Odrv4 I__2538 (
            .O(N__23917),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0 ));
    LocalMux I__2537 (
            .O(N__23914),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0 ));
    InMux I__2536 (
            .O(N__23909),
            .I(N__23906));
    LocalMux I__2535 (
            .O(N__23906),
            .I(\pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO ));
    InMux I__2534 (
            .O(N__23903),
            .I(N__23890));
    InMux I__2533 (
            .O(N__23902),
            .I(N__23890));
    InMux I__2532 (
            .O(N__23901),
            .I(N__23890));
    InMux I__2531 (
            .O(N__23900),
            .I(N__23890));
    CascadeMux I__2530 (
            .O(N__23899),
            .I(N__23886));
    LocalMux I__2529 (
            .O(N__23890),
            .I(N__23881));
    InMux I__2528 (
            .O(N__23889),
            .I(N__23876));
    InMux I__2527 (
            .O(N__23886),
            .I(N__23873));
    InMux I__2526 (
            .O(N__23885),
            .I(N__23868));
    InMux I__2525 (
            .O(N__23884),
            .I(N__23868));
    Span4Mux_v I__2524 (
            .O(N__23881),
            .I(N__23865));
    InMux I__2523 (
            .O(N__23880),
            .I(N__23860));
    InMux I__2522 (
            .O(N__23879),
            .I(N__23860));
    LocalMux I__2521 (
            .O(N__23876),
            .I(N__23857));
    LocalMux I__2520 (
            .O(N__23873),
            .I(N__23852));
    LocalMux I__2519 (
            .O(N__23868),
            .I(N__23852));
    Span4Mux_v I__2518 (
            .O(N__23865),
            .I(N__23849));
    LocalMux I__2517 (
            .O(N__23860),
            .I(N__23844));
    Span4Mux_v I__2516 (
            .O(N__23857),
            .I(N__23844));
    Odrv4 I__2515 (
            .O(N__23852),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1 ));
    Odrv4 I__2514 (
            .O(N__23849),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1 ));
    Odrv4 I__2513 (
            .O(N__23844),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1 ));
    CascadeMux I__2512 (
            .O(N__23837),
            .I(N__23834));
    InMux I__2511 (
            .O(N__23834),
            .I(N__23831));
    LocalMux I__2510 (
            .O(N__23831),
            .I(N__23827));
    CascadeMux I__2509 (
            .O(N__23830),
            .I(N__23824));
    Span4Mux_h I__2508 (
            .O(N__23827),
            .I(N__23821));
    InMux I__2507 (
            .O(N__23824),
            .I(N__23818));
    Odrv4 I__2506 (
            .O(N__23821),
            .I(\pwm_generator_inst.un18_threshold1_22 ));
    LocalMux I__2505 (
            .O(N__23818),
            .I(\pwm_generator_inst.un18_threshold1_22 ));
    InMux I__2504 (
            .O(N__23813),
            .I(N__23810));
    LocalMux I__2503 (
            .O(N__23810),
            .I(N__23807));
    Span4Mux_h I__2502 (
            .O(N__23807),
            .I(N__23803));
    InMux I__2501 (
            .O(N__23806),
            .I(N__23800));
    Odrv4 I__2500 (
            .O(N__23803),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0 ));
    LocalMux I__2499 (
            .O(N__23800),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0 ));
    CascadeMux I__2498 (
            .O(N__23795),
            .I(N__23792));
    InMux I__2497 (
            .O(N__23792),
            .I(N__23789));
    LocalMux I__2496 (
            .O(N__23789),
            .I(\pwm_generator_inst.N_179_i ));
    InMux I__2495 (
            .O(N__23786),
            .I(N__23782));
    InMux I__2494 (
            .O(N__23785),
            .I(N__23778));
    LocalMux I__2493 (
            .O(N__23782),
            .I(N__23775));
    InMux I__2492 (
            .O(N__23781),
            .I(N__23772));
    LocalMux I__2491 (
            .O(N__23778),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv12 I__2490 (
            .O(N__23775),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2489 (
            .O(N__23772),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2488 (
            .O(N__23765),
            .I(N__23762));
    LocalMux I__2487 (
            .O(N__23762),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__2486 (
            .O(N__23759),
            .I(N__23755));
    InMux I__2485 (
            .O(N__23758),
            .I(N__23751));
    LocalMux I__2484 (
            .O(N__23755),
            .I(N__23748));
    InMux I__2483 (
            .O(N__23754),
            .I(N__23745));
    LocalMux I__2482 (
            .O(N__23751),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv12 I__2481 (
            .O(N__23748),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2480 (
            .O(N__23745),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    CascadeMux I__2479 (
            .O(N__23738),
            .I(N__23735));
    InMux I__2478 (
            .O(N__23735),
            .I(N__23732));
    LocalMux I__2477 (
            .O(N__23732),
            .I(N__23729));
    Span4Mux_h I__2476 (
            .O(N__23729),
            .I(N__23726));
    Odrv4 I__2475 (
            .O(N__23726),
            .I(\pwm_generator_inst.N_180_i ));
    InMux I__2474 (
            .O(N__23723),
            .I(N__23720));
    LocalMux I__2473 (
            .O(N__23720),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__2472 (
            .O(N__23717),
            .I(N__23714));
    InMux I__2471 (
            .O(N__23714),
            .I(N__23711));
    LocalMux I__2470 (
            .O(N__23711),
            .I(\pwm_generator_inst.N_181_i ));
    CascadeMux I__2469 (
            .O(N__23708),
            .I(N__23703));
    InMux I__2468 (
            .O(N__23707),
            .I(N__23700));
    InMux I__2467 (
            .O(N__23706),
            .I(N__23697));
    InMux I__2466 (
            .O(N__23703),
            .I(N__23694));
    LocalMux I__2465 (
            .O(N__23700),
            .I(N__23691));
    LocalMux I__2464 (
            .O(N__23697),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2463 (
            .O(N__23694),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__2462 (
            .O(N__23691),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2461 (
            .O(N__23684),
            .I(N__23681));
    LocalMux I__2460 (
            .O(N__23681),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__2459 (
            .O(N__23678),
            .I(N__23673));
    InMux I__2458 (
            .O(N__23677),
            .I(N__23670));
    InMux I__2457 (
            .O(N__23676),
            .I(N__23667));
    LocalMux I__2456 (
            .O(N__23673),
            .I(N__23664));
    LocalMux I__2455 (
            .O(N__23670),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2454 (
            .O(N__23667),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__2453 (
            .O(N__23664),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    CascadeMux I__2452 (
            .O(N__23657),
            .I(N__23654));
    InMux I__2451 (
            .O(N__23654),
            .I(N__23651));
    LocalMux I__2450 (
            .O(N__23651),
            .I(\pwm_generator_inst.N_182_i ));
    InMux I__2449 (
            .O(N__23648),
            .I(N__23645));
    LocalMux I__2448 (
            .O(N__23645),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__2447 (
            .O(N__23642),
            .I(N__23639));
    InMux I__2446 (
            .O(N__23639),
            .I(N__23636));
    LocalMux I__2445 (
            .O(N__23636),
            .I(\pwm_generator_inst.N_183_i ));
    InMux I__2444 (
            .O(N__23633),
            .I(N__23628));
    InMux I__2443 (
            .O(N__23632),
            .I(N__23625));
    InMux I__2442 (
            .O(N__23631),
            .I(N__23622));
    LocalMux I__2441 (
            .O(N__23628),
            .I(N__23619));
    LocalMux I__2440 (
            .O(N__23625),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2439 (
            .O(N__23622),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__2438 (
            .O(N__23619),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2437 (
            .O(N__23612),
            .I(N__23609));
    LocalMux I__2436 (
            .O(N__23609),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__2435 (
            .O(N__23606),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2434 (
            .O(N__23603),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2433 (
            .O(N__23600),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2432 (
            .O(N__23597),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2431 (
            .O(N__23594),
            .I(bfn_3_13_0_));
    InMux I__2430 (
            .O(N__23591),
            .I(N__23573));
    InMux I__2429 (
            .O(N__23590),
            .I(N__23573));
    InMux I__2428 (
            .O(N__23589),
            .I(N__23573));
    InMux I__2427 (
            .O(N__23588),
            .I(N__23573));
    InMux I__2426 (
            .O(N__23587),
            .I(N__23568));
    InMux I__2425 (
            .O(N__23586),
            .I(N__23568));
    InMux I__2424 (
            .O(N__23585),
            .I(N__23559));
    InMux I__2423 (
            .O(N__23584),
            .I(N__23559));
    InMux I__2422 (
            .O(N__23583),
            .I(N__23559));
    InMux I__2421 (
            .O(N__23582),
            .I(N__23559));
    LocalMux I__2420 (
            .O(N__23573),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2419 (
            .O(N__23568),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2418 (
            .O(N__23559),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__2417 (
            .O(N__23552),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__2416 (
            .O(N__23549),
            .I(N__23546));
    LocalMux I__2415 (
            .O(N__23546),
            .I(\pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO ));
    InMux I__2414 (
            .O(N__23543),
            .I(N__23540));
    LocalMux I__2413 (
            .O(N__23540),
            .I(N__23537));
    Span4Mux_h I__2412 (
            .O(N__23537),
            .I(N__23533));
    InMux I__2411 (
            .O(N__23536),
            .I(N__23530));
    Odrv4 I__2410 (
            .O(N__23533),
            .I(\pwm_generator_inst.un18_threshold1_19 ));
    LocalMux I__2409 (
            .O(N__23530),
            .I(\pwm_generator_inst.un18_threshold1_19 ));
    CascadeMux I__2408 (
            .O(N__23525),
            .I(N__23522));
    InMux I__2407 (
            .O(N__23522),
            .I(N__23516));
    InMux I__2406 (
            .O(N__23521),
            .I(N__23516));
    LocalMux I__2405 (
            .O(N__23516),
            .I(N__23513));
    Span4Mux_v I__2404 (
            .O(N__23513),
            .I(N__23510));
    Odrv4 I__2403 (
            .O(N__23510),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0 ));
    InMux I__2402 (
            .O(N__23507),
            .I(N__23504));
    LocalMux I__2401 (
            .O(N__23504),
            .I(N__23501));
    Span4Mux_s3_h I__2400 (
            .O(N__23501),
            .I(N__23498));
    Odrv4 I__2399 (
            .O(N__23498),
            .I(\pwm_generator_inst.un18_threshold_1_axb_19 ));
    InMux I__2398 (
            .O(N__23495),
            .I(N__23489));
    InMux I__2397 (
            .O(N__23494),
            .I(N__23486));
    CascadeMux I__2396 (
            .O(N__23493),
            .I(N__23482));
    CascadeMux I__2395 (
            .O(N__23492),
            .I(N__23478));
    LocalMux I__2394 (
            .O(N__23489),
            .I(N__23474));
    LocalMux I__2393 (
            .O(N__23486),
            .I(N__23471));
    InMux I__2392 (
            .O(N__23485),
            .I(N__23460));
    InMux I__2391 (
            .O(N__23482),
            .I(N__23460));
    InMux I__2390 (
            .O(N__23481),
            .I(N__23460));
    InMux I__2389 (
            .O(N__23478),
            .I(N__23460));
    InMux I__2388 (
            .O(N__23477),
            .I(N__23460));
    Span4Mux_h I__2387 (
            .O(N__23474),
            .I(N__23457));
    Span12Mux_h I__2386 (
            .O(N__23471),
            .I(N__23454));
    LocalMux I__2385 (
            .O(N__23460),
            .I(N__23451));
    Span4Mux_v I__2384 (
            .O(N__23457),
            .I(N__23448));
    Span12Mux_v I__2383 (
            .O(N__23454),
            .I(N__23445));
    Span12Mux_h I__2382 (
            .O(N__23451),
            .I(N__23442));
    Span4Mux_v I__2381 (
            .O(N__23448),
            .I(N__23439));
    Odrv12 I__2380 (
            .O(N__23445),
            .I(\pwm_generator_inst.un5_threshold_1_26 ));
    Odrv12 I__2379 (
            .O(N__23442),
            .I(\pwm_generator_inst.un5_threshold_1_26 ));
    Odrv4 I__2378 (
            .O(N__23439),
            .I(\pwm_generator_inst.un5_threshold_1_26 ));
    InMux I__2377 (
            .O(N__23432),
            .I(N__23429));
    LocalMux I__2376 (
            .O(N__23429),
            .I(N__23426));
    Span4Mux_h I__2375 (
            .O(N__23426),
            .I(N__23423));
    Span4Mux_v I__2374 (
            .O(N__23423),
            .I(N__23420));
    Odrv4 I__2373 (
            .O(N__23420),
            .I(\pwm_generator_inst.un5_threshold_2_1_16 ));
    InMux I__2372 (
            .O(N__23417),
            .I(N__23414));
    LocalMux I__2371 (
            .O(N__23414),
            .I(N__23411));
    Span4Mux_v I__2370 (
            .O(N__23411),
            .I(N__23408));
    Odrv4 I__2369 (
            .O(N__23408),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0 ));
    InMux I__2368 (
            .O(N__23405),
            .I(N__23402));
    LocalMux I__2367 (
            .O(N__23402),
            .I(N__23399));
    Span4Mux_v I__2366 (
            .O(N__23399),
            .I(N__23395));
    InMux I__2365 (
            .O(N__23398),
            .I(N__23392));
    Odrv4 I__2364 (
            .O(N__23395),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0 ));
    LocalMux I__2363 (
            .O(N__23392),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0 ));
    CascadeMux I__2362 (
            .O(N__23387),
            .I(\pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_ ));
    InMux I__2361 (
            .O(N__23384),
            .I(N__23381));
    LocalMux I__2360 (
            .O(N__23381),
            .I(N__23377));
    InMux I__2359 (
            .O(N__23380),
            .I(N__23374));
    Span4Mux_v I__2358 (
            .O(N__23377),
            .I(N__23371));
    LocalMux I__2357 (
            .O(N__23374),
            .I(N__23368));
    Span4Mux_v I__2356 (
            .O(N__23371),
            .I(N__23365));
    Span4Mux_h I__2355 (
            .O(N__23368),
            .I(N__23362));
    Odrv4 I__2354 (
            .O(N__23365),
            .I(\pwm_generator_inst.un5_threshold_2_1_15 ));
    Odrv4 I__2353 (
            .O(N__23362),
            .I(\pwm_generator_inst.un5_threshold_2_1_15 ));
    InMux I__2352 (
            .O(N__23357),
            .I(N__23354));
    LocalMux I__2351 (
            .O(N__23354),
            .I(N__23351));
    Odrv4 I__2350 (
            .O(N__23351),
            .I(\pwm_generator_inst.un5_threshold_add_1_axb_16 ));
    InMux I__2349 (
            .O(N__23348),
            .I(N__23345));
    LocalMux I__2348 (
            .O(N__23345),
            .I(N__23341));
    InMux I__2347 (
            .O(N__23344),
            .I(N__23338));
    Odrv4 I__2346 (
            .O(N__23341),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0 ));
    LocalMux I__2345 (
            .O(N__23338),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0 ));
    InMux I__2344 (
            .O(N__23333),
            .I(N__23330));
    LocalMux I__2343 (
            .O(N__23330),
            .I(\pwm_generator_inst.un18_threshold_1_axb_25 ));
    InMux I__2342 (
            .O(N__23327),
            .I(N__23324));
    LocalMux I__2341 (
            .O(N__23324),
            .I(N__23321));
    Odrv4 I__2340 (
            .O(N__23321),
            .I(un8_start_stop));
    InMux I__2339 (
            .O(N__23318),
            .I(N__23315));
    LocalMux I__2338 (
            .O(N__23315),
            .I(N__23312));
    Glb2LocalMux I__2337 (
            .O(N__23312),
            .I(N__23309));
    GlobalMux I__2336 (
            .O(N__23309),
            .I(clk_12mhz));
    IoInMux I__2335 (
            .O(N__23306),
            .I(N__23303));
    LocalMux I__2334 (
            .O(N__23303),
            .I(N__23300));
    Span4Mux_s0_v I__2333 (
            .O(N__23300),
            .I(N__23297));
    Span4Mux_h I__2332 (
            .O(N__23297),
            .I(N__23294));
    Odrv4 I__2331 (
            .O(N__23294),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2330 (
            .O(N__23291),
            .I(bfn_3_12_0_));
    InMux I__2329 (
            .O(N__23288),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2328 (
            .O(N__23285),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__2327 (
            .O(N__23282),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__2326 (
            .O(N__23279),
            .I(bfn_2_16_0_));
    InMux I__2325 (
            .O(N__23276),
            .I(\pwm_generator_inst.un22_threshold_1_cry_8 ));
    InMux I__2324 (
            .O(N__23273),
            .I(N__23270));
    LocalMux I__2323 (
            .O(N__23270),
            .I(\pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO ));
    CascadeMux I__2322 (
            .O(N__23267),
            .I(N__23264));
    InMux I__2321 (
            .O(N__23264),
            .I(N__23260));
    InMux I__2320 (
            .O(N__23263),
            .I(N__23257));
    LocalMux I__2319 (
            .O(N__23260),
            .I(\pwm_generator_inst.un18_threshold1_25 ));
    LocalMux I__2318 (
            .O(N__23257),
            .I(\pwm_generator_inst.un18_threshold1_25 ));
    InMux I__2317 (
            .O(N__23252),
            .I(N__23249));
    LocalMux I__2316 (
            .O(N__23249),
            .I(\pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO ));
    InMux I__2315 (
            .O(N__23246),
            .I(N__23242));
    InMux I__2314 (
            .O(N__23245),
            .I(N__23239));
    LocalMux I__2313 (
            .O(N__23242),
            .I(\pwm_generator_inst.un22_threshold_1 ));
    LocalMux I__2312 (
            .O(N__23239),
            .I(\pwm_generator_inst.un22_threshold_1 ));
    InMux I__2311 (
            .O(N__23234),
            .I(N__23230));
    InMux I__2310 (
            .O(N__23233),
            .I(N__23227));
    LocalMux I__2309 (
            .O(N__23230),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0 ));
    LocalMux I__2308 (
            .O(N__23227),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0 ));
    InMux I__2307 (
            .O(N__23222),
            .I(N__23219));
    LocalMux I__2306 (
            .O(N__23219),
            .I(N__23216));
    Odrv4 I__2305 (
            .O(N__23216),
            .I(\pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO ));
    CascadeMux I__2304 (
            .O(N__23213),
            .I(N__23210));
    InMux I__2303 (
            .O(N__23210),
            .I(N__23207));
    LocalMux I__2302 (
            .O(N__23207),
            .I(N__23203));
    InMux I__2301 (
            .O(N__23206),
            .I(N__23200));
    Odrv4 I__2300 (
            .O(N__23203),
            .I(\pwm_generator_inst.un18_threshold1_23 ));
    LocalMux I__2299 (
            .O(N__23200),
            .I(\pwm_generator_inst.un18_threshold1_23 ));
    InMux I__2298 (
            .O(N__23195),
            .I(N__23189));
    InMux I__2297 (
            .O(N__23194),
            .I(N__23189));
    LocalMux I__2296 (
            .O(N__23189),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0 ));
    InMux I__2295 (
            .O(N__23186),
            .I(N__23183));
    LocalMux I__2294 (
            .O(N__23183),
            .I(N__23180));
    Odrv4 I__2293 (
            .O(N__23180),
            .I(\pwm_generator_inst.un18_threshold_1_axb_23 ));
    CascadeMux I__2292 (
            .O(N__23177),
            .I(N__23173));
    InMux I__2291 (
            .O(N__23176),
            .I(N__23170));
    InMux I__2290 (
            .O(N__23173),
            .I(N__23167));
    LocalMux I__2289 (
            .O(N__23170),
            .I(\pwm_generator_inst.un18_threshold1_24 ));
    LocalMux I__2288 (
            .O(N__23167),
            .I(\pwm_generator_inst.un18_threshold1_24 ));
    CascadeMux I__2287 (
            .O(N__23162),
            .I(N__23159));
    InMux I__2286 (
            .O(N__23159),
            .I(N__23156));
    LocalMux I__2285 (
            .O(N__23156),
            .I(N__23153));
    Odrv4 I__2284 (
            .O(N__23153),
            .I(\pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO ));
    InMux I__2283 (
            .O(N__23150),
            .I(N__23144));
    InMux I__2282 (
            .O(N__23149),
            .I(N__23144));
    LocalMux I__2281 (
            .O(N__23144),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0 ));
    InMux I__2280 (
            .O(N__23141),
            .I(N__23138));
    LocalMux I__2279 (
            .O(N__23138),
            .I(\pwm_generator_inst.un18_threshold_1_axb_24 ));
    InMux I__2278 (
            .O(N__23135),
            .I(N__23132));
    LocalMux I__2277 (
            .O(N__23132),
            .I(\pwm_generator_inst.un1_counterlto2_0 ));
    CascadeMux I__2276 (
            .O(N__23129),
            .I(N__23126));
    InMux I__2275 (
            .O(N__23126),
            .I(N__23122));
    CascadeMux I__2274 (
            .O(N__23125),
            .I(N__23119));
    LocalMux I__2273 (
            .O(N__23122),
            .I(N__23116));
    InMux I__2272 (
            .O(N__23119),
            .I(N__23113));
    Odrv4 I__2271 (
            .O(N__23116),
            .I(\pwm_generator_inst.un18_threshold1_18 ));
    LocalMux I__2270 (
            .O(N__23113),
            .I(\pwm_generator_inst.un18_threshold1_18 ));
    InMux I__2269 (
            .O(N__23108),
            .I(N__23105));
    LocalMux I__2268 (
            .O(N__23105),
            .I(N__23102));
    Odrv4 I__2267 (
            .O(N__23102),
            .I(\pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO ));
    InMux I__2266 (
            .O(N__23099),
            .I(\pwm_generator_inst.un22_threshold_1_cry_0 ));
    InMux I__2265 (
            .O(N__23096),
            .I(\pwm_generator_inst.un22_threshold_1_cry_1 ));
    InMux I__2264 (
            .O(N__23093),
            .I(\pwm_generator_inst.un22_threshold_1_cry_2 ));
    InMux I__2263 (
            .O(N__23090),
            .I(\pwm_generator_inst.un22_threshold_1_cry_3 ));
    InMux I__2262 (
            .O(N__23087),
            .I(\pwm_generator_inst.un22_threshold_1_cry_4 ));
    InMux I__2261 (
            .O(N__23084),
            .I(\pwm_generator_inst.un22_threshold_1_cry_5 ));
    InMux I__2260 (
            .O(N__23081),
            .I(\pwm_generator_inst.un22_threshold_1_cry_6 ));
    InMux I__2259 (
            .O(N__23078),
            .I(\pwm_generator_inst.un3_threshold_cry_16 ));
    InMux I__2258 (
            .O(N__23075),
            .I(N__23072));
    LocalMux I__2257 (
            .O(N__23072),
            .I(N__23069));
    Span4Mux_s1_h I__2256 (
            .O(N__23069),
            .I(N__23066));
    Odrv4 I__2255 (
            .O(N__23066),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0 ));
    InMux I__2254 (
            .O(N__23063),
            .I(\pwm_generator_inst.un3_threshold_cry_17 ));
    InMux I__2253 (
            .O(N__23060),
            .I(\pwm_generator_inst.un3_threshold_cry_18 ));
    InMux I__2252 (
            .O(N__23057),
            .I(N__23054));
    LocalMux I__2251 (
            .O(N__23054),
            .I(N__23051));
    Span4Mux_v I__2250 (
            .O(N__23051),
            .I(N__23048));
    Odrv4 I__2249 (
            .O(N__23048),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__2248 (
            .O(N__23045),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    CascadeMux I__2247 (
            .O(N__23042),
            .I(N__23039));
    InMux I__2246 (
            .O(N__23039),
            .I(N__23036));
    LocalMux I__2245 (
            .O(N__23036),
            .I(N__23033));
    Span4Mux_v I__2244 (
            .O(N__23033),
            .I(N__23030));
    Odrv4 I__2243 (
            .O(N__23030),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0 ));
    InMux I__2242 (
            .O(N__23027),
            .I(N__23024));
    LocalMux I__2241 (
            .O(N__23024),
            .I(N_112_i_i));
    InMux I__2240 (
            .O(N__23021),
            .I(N__23018));
    LocalMux I__2239 (
            .O(N__23018),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    CascadeMux I__2238 (
            .O(N__23015),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__2237 (
            .O(N__23012),
            .I(N__23009));
    LocalMux I__2236 (
            .O(N__23009),
            .I(N__23006));
    Span4Mux_h I__2235 (
            .O(N__23006),
            .I(N__23002));
    InMux I__2234 (
            .O(N__23005),
            .I(N__22999));
    Odrv4 I__2233 (
            .O(N__23002),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0 ));
    LocalMux I__2232 (
            .O(N__22999),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0 ));
    InMux I__2231 (
            .O(N__22994),
            .I(N__22991));
    LocalMux I__2230 (
            .O(N__22991),
            .I(N__22988));
    Span4Mux_v I__2229 (
            .O(N__22988),
            .I(N__22985));
    Odrv4 I__2228 (
            .O(N__22985),
            .I(\pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8 ));
    InMux I__2227 (
            .O(N__22982),
            .I(\pwm_generator_inst.un3_threshold_cry_8 ));
    InMux I__2226 (
            .O(N__22979),
            .I(N__22976));
    LocalMux I__2225 (
            .O(N__22976),
            .I(N__22973));
    Span4Mux_v I__2224 (
            .O(N__22973),
            .I(N__22970));
    Odrv4 I__2223 (
            .O(N__22970),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8 ));
    InMux I__2222 (
            .O(N__22967),
            .I(\pwm_generator_inst.un3_threshold_cry_9 ));
    InMux I__2221 (
            .O(N__22964),
            .I(N__22961));
    LocalMux I__2220 (
            .O(N__22961),
            .I(N__22958));
    Span4Mux_v I__2219 (
            .O(N__22958),
            .I(N__22955));
    Odrv4 I__2218 (
            .O(N__22955),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7 ));
    InMux I__2217 (
            .O(N__22952),
            .I(\pwm_generator_inst.un3_threshold_cry_10 ));
    InMux I__2216 (
            .O(N__22949),
            .I(N__22946));
    LocalMux I__2215 (
            .O(N__22946),
            .I(N__22943));
    Span4Mux_v I__2214 (
            .O(N__22943),
            .I(N__22940));
    Odrv4 I__2213 (
            .O(N__22940),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7 ));
    InMux I__2212 (
            .O(N__22937),
            .I(\pwm_generator_inst.un3_threshold_cry_11 ));
    InMux I__2211 (
            .O(N__22934),
            .I(N__22931));
    LocalMux I__2210 (
            .O(N__22931),
            .I(N__22928));
    Span4Mux_v I__2209 (
            .O(N__22928),
            .I(N__22925));
    Odrv4 I__2208 (
            .O(N__22925),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7 ));
    InMux I__2207 (
            .O(N__22922),
            .I(\pwm_generator_inst.un3_threshold_cry_12 ));
    InMux I__2206 (
            .O(N__22919),
            .I(N__22916));
    LocalMux I__2205 (
            .O(N__22916),
            .I(N__22913));
    Span4Mux_v I__2204 (
            .O(N__22913),
            .I(N__22910));
    Odrv4 I__2203 (
            .O(N__22910),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7 ));
    InMux I__2202 (
            .O(N__22907),
            .I(\pwm_generator_inst.un3_threshold_cry_13 ));
    InMux I__2201 (
            .O(N__22904),
            .I(N__22901));
    LocalMux I__2200 (
            .O(N__22901),
            .I(N__22898));
    Span4Mux_v I__2199 (
            .O(N__22898),
            .I(N__22895));
    Odrv4 I__2198 (
            .O(N__22895),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7 ));
    InMux I__2197 (
            .O(N__22892),
            .I(\pwm_generator_inst.un3_threshold_cry_14 ));
    InMux I__2196 (
            .O(N__22889),
            .I(N__22886));
    LocalMux I__2195 (
            .O(N__22886),
            .I(N__22883));
    Span4Mux_v I__2194 (
            .O(N__22883),
            .I(N__22880));
    Odrv4 I__2193 (
            .O(N__22880),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7 ));
    InMux I__2192 (
            .O(N__22877),
            .I(bfn_1_22_0_));
    InMux I__2191 (
            .O(N__22874),
            .I(N__22871));
    LocalMux I__2190 (
            .O(N__22871),
            .I(N__22868));
    Span4Mux_v I__2189 (
            .O(N__22868),
            .I(N__22865));
    Odrv4 I__2188 (
            .O(N__22865),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7 ));
    InMux I__2187 (
            .O(N__22862),
            .I(N__22859));
    LocalMux I__2186 (
            .O(N__22859),
            .I(N__22856));
    Span12Mux_v I__2185 (
            .O(N__22856),
            .I(N__22853));
    Span12Mux_h I__2184 (
            .O(N__22853),
            .I(N__22850));
    Span12Mux_h I__2183 (
            .O(N__22850),
            .I(N__22847));
    Odrv12 I__2182 (
            .O(N__22847),
            .I(\pwm_generator_inst.O_0_8 ));
    InMux I__2181 (
            .O(N__22844),
            .I(N__22841));
    LocalMux I__2180 (
            .O(N__22841),
            .I(N__22838));
    Span4Mux_v I__2179 (
            .O(N__22838),
            .I(N__22835));
    Sp12to4 I__2178 (
            .O(N__22835),
            .I(N__22832));
    Odrv12 I__2177 (
            .O(N__22832),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0 ));
    InMux I__2176 (
            .O(N__22829),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    CascadeMux I__2175 (
            .O(N__22826),
            .I(N__22823));
    InMux I__2174 (
            .O(N__22823),
            .I(N__22820));
    LocalMux I__2173 (
            .O(N__22820),
            .I(N__22817));
    Span12Mux_v I__2172 (
            .O(N__22817),
            .I(N__22814));
    Span12Mux_h I__2171 (
            .O(N__22814),
            .I(N__22811));
    Span12Mux_h I__2170 (
            .O(N__22811),
            .I(N__22808));
    Odrv12 I__2169 (
            .O(N__22808),
            .I(\pwm_generator_inst.O_0_9 ));
    InMux I__2168 (
            .O(N__22805),
            .I(N__22802));
    LocalMux I__2167 (
            .O(N__22802),
            .I(N__22799));
    Span4Mux_v I__2166 (
            .O(N__22799),
            .I(N__22796));
    Sp12to4 I__2165 (
            .O(N__22796),
            .I(N__22793));
    Odrv12 I__2164 (
            .O(N__22793),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0 ));
    InMux I__2163 (
            .O(N__22790),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__2162 (
            .O(N__22787),
            .I(N__22784));
    LocalMux I__2161 (
            .O(N__22784),
            .I(N__22781));
    Span12Mux_v I__2160 (
            .O(N__22781),
            .I(N__22778));
    Span12Mux_h I__2159 (
            .O(N__22778),
            .I(N__22775));
    Span12Mux_h I__2158 (
            .O(N__22775),
            .I(N__22772));
    Odrv12 I__2157 (
            .O(N__22772),
            .I(\pwm_generator_inst.O_0_10 ));
    InMux I__2156 (
            .O(N__22769),
            .I(N__22766));
    LocalMux I__2155 (
            .O(N__22766),
            .I(N__22763));
    Span12Mux_s1_h I__2154 (
            .O(N__22763),
            .I(N__22760));
    Span12Mux_v I__2153 (
            .O(N__22760),
            .I(N__22757));
    Odrv12 I__2152 (
            .O(N__22757),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0 ));
    InMux I__2151 (
            .O(N__22754),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__2150 (
            .O(N__22751),
            .I(N__22748));
    LocalMux I__2149 (
            .O(N__22748),
            .I(N__22745));
    Span12Mux_v I__2148 (
            .O(N__22745),
            .I(N__22742));
    Span12Mux_h I__2147 (
            .O(N__22742),
            .I(N__22739));
    Span12Mux_h I__2146 (
            .O(N__22739),
            .I(N__22736));
    Odrv12 I__2145 (
            .O(N__22736),
            .I(\pwm_generator_inst.O_0_11 ));
    InMux I__2144 (
            .O(N__22733),
            .I(N__22730));
    LocalMux I__2143 (
            .O(N__22730),
            .I(N__22727));
    Span4Mux_v I__2142 (
            .O(N__22727),
            .I(N__22724));
    Odrv4 I__2141 (
            .O(N__22724),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0 ));
    InMux I__2140 (
            .O(N__22721),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__2139 (
            .O(N__22718),
            .I(N__22715));
    LocalMux I__2138 (
            .O(N__22715),
            .I(N__22712));
    Span12Mux_h I__2137 (
            .O(N__22712),
            .I(N__22709));
    Span12Mux_h I__2136 (
            .O(N__22709),
            .I(N__22706));
    Odrv12 I__2135 (
            .O(N__22706),
            .I(\pwm_generator_inst.O_0_12 ));
    InMux I__2134 (
            .O(N__22703),
            .I(N__22700));
    LocalMux I__2133 (
            .O(N__22700),
            .I(N__22697));
    Span4Mux_v I__2132 (
            .O(N__22697),
            .I(N__22694));
    Odrv4 I__2131 (
            .O(N__22694),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0 ));
    InMux I__2130 (
            .O(N__22691),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__2129 (
            .O(N__22688),
            .I(N__22685));
    LocalMux I__2128 (
            .O(N__22685),
            .I(N__22682));
    Span4Mux_v I__2127 (
            .O(N__22682),
            .I(N__22679));
    Sp12to4 I__2126 (
            .O(N__22679),
            .I(N__22676));
    Span12Mux_h I__2125 (
            .O(N__22676),
            .I(N__22673));
    Span12Mux_h I__2124 (
            .O(N__22673),
            .I(N__22670));
    Odrv12 I__2123 (
            .O(N__22670),
            .I(\pwm_generator_inst.O_0_13 ));
    InMux I__2122 (
            .O(N__22667),
            .I(N__22664));
    LocalMux I__2121 (
            .O(N__22664),
            .I(N__22661));
    Span4Mux_v I__2120 (
            .O(N__22661),
            .I(N__22658));
    Odrv4 I__2119 (
            .O(N__22658),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0 ));
    InMux I__2118 (
            .O(N__22655),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__2117 (
            .O(N__22652),
            .I(N__22649));
    LocalMux I__2116 (
            .O(N__22649),
            .I(N__22646));
    Span4Mux_v I__2115 (
            .O(N__22646),
            .I(N__22643));
    Sp12to4 I__2114 (
            .O(N__22643),
            .I(N__22640));
    Span12Mux_h I__2113 (
            .O(N__22640),
            .I(N__22637));
    Odrv12 I__2112 (
            .O(N__22637),
            .I(\pwm_generator_inst.O_0_14 ));
    InMux I__2111 (
            .O(N__22634),
            .I(N__22631));
    LocalMux I__2110 (
            .O(N__22631),
            .I(N__22628));
    Span4Mux_v I__2109 (
            .O(N__22628),
            .I(N__22625));
    Odrv4 I__2108 (
            .O(N__22625),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0 ));
    InMux I__2107 (
            .O(N__22622),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__2106 (
            .O(N__22619),
            .I(N__22616));
    LocalMux I__2105 (
            .O(N__22616),
            .I(N__22613));
    Span4Mux_v I__2104 (
            .O(N__22613),
            .I(N__22610));
    Odrv4 I__2103 (
            .O(N__22610),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0 ));
    InMux I__2102 (
            .O(N__22607),
            .I(bfn_1_21_0_));
    InMux I__2101 (
            .O(N__22604),
            .I(N__22601));
    LocalMux I__2100 (
            .O(N__22601),
            .I(N__22598));
    Span4Mux_v I__2099 (
            .O(N__22598),
            .I(N__22595));
    Span4Mux_v I__2098 (
            .O(N__22595),
            .I(N__22592));
    Odrv4 I__2097 (
            .O(N__22592),
            .I(\pwm_generator_inst.un5_threshold_1_25 ));
    CascadeMux I__2096 (
            .O(N__22589),
            .I(N__22586));
    InMux I__2095 (
            .O(N__22586),
            .I(N__22583));
    LocalMux I__2094 (
            .O(N__22583),
            .I(N__22580));
    Span4Mux_v I__2093 (
            .O(N__22580),
            .I(N__22577));
    Odrv4 I__2092 (
            .O(N__22577),
            .I(\pwm_generator_inst.un5_threshold_2_10 ));
    InMux I__2091 (
            .O(N__22574),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_9 ));
    CascadeMux I__2090 (
            .O(N__22571),
            .I(N__22568));
    InMux I__2089 (
            .O(N__22568),
            .I(N__22565));
    LocalMux I__2088 (
            .O(N__22565),
            .I(N__22562));
    Span4Mux_v I__2087 (
            .O(N__22562),
            .I(N__22559));
    Odrv4 I__2086 (
            .O(N__22559),
            .I(\pwm_generator_inst.un5_threshold_2_11 ));
    InMux I__2085 (
            .O(N__22556),
            .I(N__22553));
    LocalMux I__2084 (
            .O(N__22553),
            .I(N__22550));
    Odrv4 I__2083 (
            .O(N__22550),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0 ));
    InMux I__2082 (
            .O(N__22547),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_10 ));
    InMux I__2081 (
            .O(N__22544),
            .I(N__22541));
    LocalMux I__2080 (
            .O(N__22541),
            .I(N__22538));
    Span4Mux_v I__2079 (
            .O(N__22538),
            .I(N__22535));
    Odrv4 I__2078 (
            .O(N__22535),
            .I(\pwm_generator_inst.un5_threshold_2_12 ));
    CascadeMux I__2077 (
            .O(N__22532),
            .I(N__22529));
    InMux I__2076 (
            .O(N__22529),
            .I(N__22526));
    LocalMux I__2075 (
            .O(N__22526),
            .I(N__22523));
    Span4Mux_v I__2074 (
            .O(N__22523),
            .I(N__22520));
    Odrv4 I__2073 (
            .O(N__22520),
            .I(\pwm_generator_inst.un5_threshold_2_13 ));
    InMux I__2072 (
            .O(N__22517),
            .I(N__22514));
    LocalMux I__2071 (
            .O(N__22514),
            .I(N__22511));
    Span4Mux_v I__2070 (
            .O(N__22511),
            .I(N__22508));
    Odrv4 I__2069 (
            .O(N__22508),
            .I(\pwm_generator_inst.un5_threshold_2_14 ));
    InMux I__2068 (
            .O(N__22505),
            .I(bfn_1_19_0_));
    InMux I__2067 (
            .O(N__22502),
            .I(N__22499));
    LocalMux I__2066 (
            .O(N__22499),
            .I(N__22496));
    Span4Mux_v I__2065 (
            .O(N__22496),
            .I(N__22493));
    Odrv4 I__2064 (
            .O(N__22493),
            .I(\pwm_generator_inst.un5_threshold_2_2 ));
    CascadeMux I__2063 (
            .O(N__22490),
            .I(N__22487));
    InMux I__2062 (
            .O(N__22487),
            .I(N__22484));
    LocalMux I__2061 (
            .O(N__22484),
            .I(N__22481));
    Span4Mux_v I__2060 (
            .O(N__22481),
            .I(N__22478));
    Span4Mux_v I__2059 (
            .O(N__22478),
            .I(N__22475));
    Odrv4 I__2058 (
            .O(N__22475),
            .I(\pwm_generator_inst.un5_threshold_1_17 ));
    InMux I__2057 (
            .O(N__22472),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_1 ));
    InMux I__2056 (
            .O(N__22469),
            .I(N__22466));
    LocalMux I__2055 (
            .O(N__22466),
            .I(N__22463));
    Span4Mux_v I__2054 (
            .O(N__22463),
            .I(N__22460));
    Odrv4 I__2053 (
            .O(N__22460),
            .I(\pwm_generator_inst.un5_threshold_2_3 ));
    CascadeMux I__2052 (
            .O(N__22457),
            .I(N__22454));
    InMux I__2051 (
            .O(N__22454),
            .I(N__22451));
    LocalMux I__2050 (
            .O(N__22451),
            .I(N__22448));
    Span4Mux_v I__2049 (
            .O(N__22448),
            .I(N__22445));
    Span4Mux_s1_h I__2048 (
            .O(N__22445),
            .I(N__22442));
    Span4Mux_v I__2047 (
            .O(N__22442),
            .I(N__22439));
    Odrv4 I__2046 (
            .O(N__22439),
            .I(\pwm_generator_inst.un5_threshold_1_18 ));
    InMux I__2045 (
            .O(N__22436),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_2 ));
    InMux I__2044 (
            .O(N__22433),
            .I(N__22430));
    LocalMux I__2043 (
            .O(N__22430),
            .I(N__22427));
    Span4Mux_v I__2042 (
            .O(N__22427),
            .I(N__22424));
    Odrv4 I__2041 (
            .O(N__22424),
            .I(\pwm_generator_inst.un5_threshold_2_4 ));
    CascadeMux I__2040 (
            .O(N__22421),
            .I(N__22418));
    InMux I__2039 (
            .O(N__22418),
            .I(N__22415));
    LocalMux I__2038 (
            .O(N__22415),
            .I(N__22412));
    Span4Mux_v I__2037 (
            .O(N__22412),
            .I(N__22409));
    Span4Mux_v I__2036 (
            .O(N__22409),
            .I(N__22406));
    Odrv4 I__2035 (
            .O(N__22406),
            .I(\pwm_generator_inst.un5_threshold_1_19 ));
    InMux I__2034 (
            .O(N__22403),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_3 ));
    InMux I__2033 (
            .O(N__22400),
            .I(N__22397));
    LocalMux I__2032 (
            .O(N__22397),
            .I(N__22394));
    Span4Mux_v I__2031 (
            .O(N__22394),
            .I(N__22391));
    Odrv4 I__2030 (
            .O(N__22391),
            .I(\pwm_generator_inst.un5_threshold_2_5 ));
    CascadeMux I__2029 (
            .O(N__22388),
            .I(N__22385));
    InMux I__2028 (
            .O(N__22385),
            .I(N__22382));
    LocalMux I__2027 (
            .O(N__22382),
            .I(N__22379));
    Span4Mux_v I__2026 (
            .O(N__22379),
            .I(N__22376));
    Span4Mux_v I__2025 (
            .O(N__22376),
            .I(N__22373));
    Odrv4 I__2024 (
            .O(N__22373),
            .I(\pwm_generator_inst.un5_threshold_1_20 ));
    InMux I__2023 (
            .O(N__22370),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_4 ));
    InMux I__2022 (
            .O(N__22367),
            .I(N__22364));
    LocalMux I__2021 (
            .O(N__22364),
            .I(N__22361));
    Span4Mux_v I__2020 (
            .O(N__22361),
            .I(N__22358));
    Span4Mux_v I__2019 (
            .O(N__22358),
            .I(N__22355));
    Odrv4 I__2018 (
            .O(N__22355),
            .I(\pwm_generator_inst.un5_threshold_1_21 ));
    CascadeMux I__2017 (
            .O(N__22352),
            .I(N__22349));
    InMux I__2016 (
            .O(N__22349),
            .I(N__22346));
    LocalMux I__2015 (
            .O(N__22346),
            .I(N__22343));
    Span4Mux_v I__2014 (
            .O(N__22343),
            .I(N__22340));
    Odrv4 I__2013 (
            .O(N__22340),
            .I(\pwm_generator_inst.un5_threshold_2_6 ));
    InMux I__2012 (
            .O(N__22337),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_5 ));
    InMux I__2011 (
            .O(N__22334),
            .I(N__22331));
    LocalMux I__2010 (
            .O(N__22331),
            .I(N__22328));
    Span4Mux_v I__2009 (
            .O(N__22328),
            .I(N__22325));
    Span4Mux_v I__2008 (
            .O(N__22325),
            .I(N__22322));
    Odrv4 I__2007 (
            .O(N__22322),
            .I(\pwm_generator_inst.un5_threshold_1_22 ));
    CascadeMux I__2006 (
            .O(N__22319),
            .I(N__22316));
    InMux I__2005 (
            .O(N__22316),
            .I(N__22313));
    LocalMux I__2004 (
            .O(N__22313),
            .I(N__22310));
    Span4Mux_v I__2003 (
            .O(N__22310),
            .I(N__22307));
    Odrv4 I__2002 (
            .O(N__22307),
            .I(\pwm_generator_inst.un5_threshold_2_7 ));
    InMux I__2001 (
            .O(N__22304),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_6 ));
    InMux I__2000 (
            .O(N__22301),
            .I(N__22298));
    LocalMux I__1999 (
            .O(N__22298),
            .I(N__22295));
    Span4Mux_v I__1998 (
            .O(N__22295),
            .I(N__22292));
    Span4Mux_v I__1997 (
            .O(N__22292),
            .I(N__22289));
    Odrv4 I__1996 (
            .O(N__22289),
            .I(\pwm_generator_inst.un5_threshold_1_23 ));
    CascadeMux I__1995 (
            .O(N__22286),
            .I(N__22283));
    InMux I__1994 (
            .O(N__22283),
            .I(N__22280));
    LocalMux I__1993 (
            .O(N__22280),
            .I(N__22277));
    Span4Mux_v I__1992 (
            .O(N__22277),
            .I(N__22274));
    Odrv4 I__1991 (
            .O(N__22274),
            .I(\pwm_generator_inst.un5_threshold_2_8 ));
    InMux I__1990 (
            .O(N__22271),
            .I(bfn_1_18_0_));
    InMux I__1989 (
            .O(N__22268),
            .I(N__22265));
    LocalMux I__1988 (
            .O(N__22265),
            .I(N__22262));
    Span4Mux_v I__1987 (
            .O(N__22262),
            .I(N__22259));
    Span4Mux_v I__1986 (
            .O(N__22259),
            .I(N__22256));
    Odrv4 I__1985 (
            .O(N__22256),
            .I(\pwm_generator_inst.un5_threshold_1_24 ));
    CascadeMux I__1984 (
            .O(N__22253),
            .I(N__22250));
    InMux I__1983 (
            .O(N__22250),
            .I(N__22247));
    LocalMux I__1982 (
            .O(N__22247),
            .I(N__22244));
    Span4Mux_v I__1981 (
            .O(N__22244),
            .I(N__22241));
    Odrv4 I__1980 (
            .O(N__22241),
            .I(\pwm_generator_inst.un5_threshold_2_9 ));
    InMux I__1979 (
            .O(N__22238),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_8 ));
    InMux I__1978 (
            .O(N__22235),
            .I(\pwm_generator_inst.un18_threshold_1_cry_24 ));
    InMux I__1977 (
            .O(N__22232),
            .I(\pwm_generator_inst.un18_threshold_1_cry_25 ));
    InMux I__1976 (
            .O(N__22229),
            .I(N__22226));
    LocalMux I__1975 (
            .O(N__22226),
            .I(\pwm_generator_inst.un18_threshold_1_axb_20 ));
    InMux I__1974 (
            .O(N__22223),
            .I(N__22220));
    LocalMux I__1973 (
            .O(N__22220),
            .I(\pwm_generator_inst.un18_threshold_1_axb_17 ));
    InMux I__1972 (
            .O(N__22217),
            .I(N__22214));
    LocalMux I__1971 (
            .O(N__22214),
            .I(\pwm_generator_inst.un18_threshold_1_axb_18 ));
    InMux I__1970 (
            .O(N__22211),
            .I(N__22208));
    LocalMux I__1969 (
            .O(N__22208),
            .I(\pwm_generator_inst.un18_threshold_1_axb_22 ));
    InMux I__1968 (
            .O(N__22205),
            .I(N__22202));
    LocalMux I__1967 (
            .O(N__22202),
            .I(\pwm_generator_inst.un18_threshold_1_axb_21 ));
    InMux I__1966 (
            .O(N__22199),
            .I(N__22196));
    LocalMux I__1965 (
            .O(N__22196),
            .I(N__22193));
    Span4Mux_v I__1964 (
            .O(N__22193),
            .I(N__22190));
    Odrv4 I__1963 (
            .O(N__22190),
            .I(\pwm_generator_inst.un5_threshold_2_0 ));
    CascadeMux I__1962 (
            .O(N__22187),
            .I(N__22184));
    InMux I__1961 (
            .O(N__22184),
            .I(N__22181));
    LocalMux I__1960 (
            .O(N__22181),
            .I(N__22178));
    Span12Mux_v I__1959 (
            .O(N__22178),
            .I(N__22175));
    Odrv12 I__1958 (
            .O(N__22175),
            .I(\pwm_generator_inst.un5_threshold_1_15 ));
    InMux I__1957 (
            .O(N__22172),
            .I(N__22169));
    LocalMux I__1956 (
            .O(N__22169),
            .I(N__22166));
    Odrv4 I__1955 (
            .O(N__22166),
            .I(\pwm_generator_inst.un18_threshold_1_axb_15 ));
    InMux I__1954 (
            .O(N__22163),
            .I(N__22160));
    LocalMux I__1953 (
            .O(N__22160),
            .I(N__22157));
    Span4Mux_v I__1952 (
            .O(N__22157),
            .I(N__22154));
    Odrv4 I__1951 (
            .O(N__22154),
            .I(\pwm_generator_inst.un5_threshold_2_1 ));
    CascadeMux I__1950 (
            .O(N__22151),
            .I(N__22148));
    InMux I__1949 (
            .O(N__22148),
            .I(N__22145));
    LocalMux I__1948 (
            .O(N__22145),
            .I(N__22142));
    Span4Mux_v I__1947 (
            .O(N__22142),
            .I(N__22139));
    Span4Mux_v I__1946 (
            .O(N__22139),
            .I(N__22136));
    Odrv4 I__1945 (
            .O(N__22136),
            .I(\pwm_generator_inst.un5_threshold_1_16 ));
    InMux I__1944 (
            .O(N__22133),
            .I(N__22130));
    LocalMux I__1943 (
            .O(N__22130),
            .I(N__22127));
    Odrv4 I__1942 (
            .O(N__22127),
            .I(\pwm_generator_inst.un18_threshold_1_axb_16 ));
    InMux I__1941 (
            .O(N__22124),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_0 ));
    InMux I__1940 (
            .O(N__22121),
            .I(\pwm_generator_inst.un18_threshold_1_cry_16 ));
    InMux I__1939 (
            .O(N__22118),
            .I(\pwm_generator_inst.un18_threshold_1_cry_17 ));
    InMux I__1938 (
            .O(N__22115),
            .I(\pwm_generator_inst.un18_threshold_1_cry_18 ));
    InMux I__1937 (
            .O(N__22112),
            .I(\pwm_generator_inst.un18_threshold_1_cry_19 ));
    InMux I__1936 (
            .O(N__22109),
            .I(\pwm_generator_inst.un18_threshold_1_cry_20 ));
    InMux I__1935 (
            .O(N__22106),
            .I(\pwm_generator_inst.un18_threshold_1_cry_21 ));
    InMux I__1934 (
            .O(N__22103),
            .I(\pwm_generator_inst.un18_threshold_1_cry_22 ));
    InMux I__1933 (
            .O(N__22100),
            .I(bfn_1_16_0_));
    InMux I__1932 (
            .O(N__22097),
            .I(N__22094));
    LocalMux I__1931 (
            .O(N__22094),
            .I(N__22091));
    Span12Mux_h I__1930 (
            .O(N__22091),
            .I(N__22088));
    Odrv12 I__1929 (
            .O(N__22088),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1928 (
            .O(N__22085),
            .I(N__22082));
    LocalMux I__1927 (
            .O(N__22082),
            .I(\pwm_generator_inst.un18_threshold_1_axb_8 ));
    InMux I__1926 (
            .O(N__22079),
            .I(N__22076));
    LocalMux I__1925 (
            .O(N__22076),
            .I(N__22073));
    Span4Mux_v I__1924 (
            .O(N__22073),
            .I(N__22070));
    Span4Mux_v I__1923 (
            .O(N__22070),
            .I(N__22067));
    Odrv4 I__1922 (
            .O(N__22067),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1921 (
            .O(N__22064),
            .I(N__22061));
    LocalMux I__1920 (
            .O(N__22061),
            .I(\pwm_generator_inst.un18_threshold_1_axb_9 ));
    InMux I__1919 (
            .O(N__22058),
            .I(N__22055));
    LocalMux I__1918 (
            .O(N__22055),
            .I(N__22052));
    Span4Mux_v I__1917 (
            .O(N__22052),
            .I(N__22049));
    Span4Mux_v I__1916 (
            .O(N__22049),
            .I(N__22046));
    Odrv4 I__1915 (
            .O(N__22046),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1914 (
            .O(N__22043),
            .I(N__22040));
    LocalMux I__1913 (
            .O(N__22040),
            .I(\pwm_generator_inst.un18_threshold_1_axb_10 ));
    InMux I__1912 (
            .O(N__22037),
            .I(N__22034));
    LocalMux I__1911 (
            .O(N__22034),
            .I(N__22031));
    Span4Mux_v I__1910 (
            .O(N__22031),
            .I(N__22028));
    Span4Mux_v I__1909 (
            .O(N__22028),
            .I(N__22025));
    Odrv4 I__1908 (
            .O(N__22025),
            .I(\pwm_generator_inst.O_11 ));
    InMux I__1907 (
            .O(N__22022),
            .I(N__22019));
    LocalMux I__1906 (
            .O(N__22019),
            .I(\pwm_generator_inst.un18_threshold_1_axb_11 ));
    InMux I__1905 (
            .O(N__22016),
            .I(N__22013));
    LocalMux I__1904 (
            .O(N__22013),
            .I(N__22010));
    Span4Mux_v I__1903 (
            .O(N__22010),
            .I(N__22007));
    Span4Mux_v I__1902 (
            .O(N__22007),
            .I(N__22004));
    Odrv4 I__1901 (
            .O(N__22004),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1900 (
            .O(N__22001),
            .I(N__21998));
    LocalMux I__1899 (
            .O(N__21998),
            .I(\pwm_generator_inst.un18_threshold_1_axb_12 ));
    InMux I__1898 (
            .O(N__21995),
            .I(N__21992));
    LocalMux I__1897 (
            .O(N__21992),
            .I(N__21989));
    Span4Mux_v I__1896 (
            .O(N__21989),
            .I(N__21986));
    Span4Mux_v I__1895 (
            .O(N__21986),
            .I(N__21983));
    Odrv4 I__1894 (
            .O(N__21983),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1893 (
            .O(N__21980),
            .I(N__21977));
    LocalMux I__1892 (
            .O(N__21977),
            .I(\pwm_generator_inst.un18_threshold_1_axb_13 ));
    InMux I__1891 (
            .O(N__21974),
            .I(N__21971));
    LocalMux I__1890 (
            .O(N__21971),
            .I(N__21968));
    Span4Mux_v I__1889 (
            .O(N__21968),
            .I(N__21965));
    Span4Mux_v I__1888 (
            .O(N__21965),
            .I(N__21962));
    Odrv4 I__1887 (
            .O(N__21962),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1886 (
            .O(N__21959),
            .I(N__21956));
    LocalMux I__1885 (
            .O(N__21956),
            .I(\pwm_generator_inst.un18_threshold_1_axb_14 ));
    InMux I__1884 (
            .O(N__21953),
            .I(N__21950));
    LocalMux I__1883 (
            .O(N__21950),
            .I(N__21947));
    Span4Mux_v I__1882 (
            .O(N__21947),
            .I(N__21944));
    Span4Mux_v I__1881 (
            .O(N__21944),
            .I(N__21941));
    Odrv4 I__1880 (
            .O(N__21941),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1879 (
            .O(N__21938),
            .I(N__21935));
    LocalMux I__1878 (
            .O(N__21935),
            .I(\pwm_generator_inst.un18_threshold_1_axb_1 ));
    InMux I__1877 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__1876 (
            .O(N__21929),
            .I(N__21926));
    Span4Mux_v I__1875 (
            .O(N__21926),
            .I(N__21923));
    Span4Mux_v I__1874 (
            .O(N__21923),
            .I(N__21920));
    Odrv4 I__1873 (
            .O(N__21920),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1872 (
            .O(N__21917),
            .I(N__21914));
    LocalMux I__1871 (
            .O(N__21914),
            .I(\pwm_generator_inst.un18_threshold_1_axb_2 ));
    InMux I__1870 (
            .O(N__21911),
            .I(N__21908));
    LocalMux I__1869 (
            .O(N__21908),
            .I(N__21905));
    Span4Mux_v I__1868 (
            .O(N__21905),
            .I(N__21902));
    Span4Mux_v I__1867 (
            .O(N__21902),
            .I(N__21899));
    Odrv4 I__1866 (
            .O(N__21899),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1865 (
            .O(N__21896),
            .I(N__21893));
    LocalMux I__1864 (
            .O(N__21893),
            .I(\pwm_generator_inst.un18_threshold_1_axb_3 ));
    InMux I__1863 (
            .O(N__21890),
            .I(N__21887));
    LocalMux I__1862 (
            .O(N__21887),
            .I(N__21884));
    Span4Mux_v I__1861 (
            .O(N__21884),
            .I(N__21881));
    Span4Mux_v I__1860 (
            .O(N__21881),
            .I(N__21878));
    Odrv4 I__1859 (
            .O(N__21878),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1858 (
            .O(N__21875),
            .I(N__21872));
    LocalMux I__1857 (
            .O(N__21872),
            .I(\pwm_generator_inst.un18_threshold_1_axb_4 ));
    InMux I__1856 (
            .O(N__21869),
            .I(N__21866));
    LocalMux I__1855 (
            .O(N__21866),
            .I(N__21863));
    Span4Mux_v I__1854 (
            .O(N__21863),
            .I(N__21860));
    Span4Mux_v I__1853 (
            .O(N__21860),
            .I(N__21857));
    Odrv4 I__1852 (
            .O(N__21857),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1851 (
            .O(N__21854),
            .I(N__21851));
    LocalMux I__1850 (
            .O(N__21851),
            .I(\pwm_generator_inst.un18_threshold_1_axb_5 ));
    InMux I__1849 (
            .O(N__21848),
            .I(N__21845));
    LocalMux I__1848 (
            .O(N__21845),
            .I(N__21842));
    Span4Mux_v I__1847 (
            .O(N__21842),
            .I(N__21839));
    Span4Mux_v I__1846 (
            .O(N__21839),
            .I(N__21836));
    Odrv4 I__1845 (
            .O(N__21836),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1844 (
            .O(N__21833),
            .I(N__21830));
    LocalMux I__1843 (
            .O(N__21830),
            .I(\pwm_generator_inst.un18_threshold_1_axb_6 ));
    InMux I__1842 (
            .O(N__21827),
            .I(N__21824));
    LocalMux I__1841 (
            .O(N__21824),
            .I(N__21821));
    Span12Mux_v I__1840 (
            .O(N__21821),
            .I(N__21818));
    Odrv12 I__1839 (
            .O(N__21818),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1838 (
            .O(N__21815),
            .I(N__21812));
    LocalMux I__1837 (
            .O(N__21812),
            .I(\pwm_generator_inst.un18_threshold_1_axb_7 ));
    InMux I__1836 (
            .O(N__21809),
            .I(N__21806));
    LocalMux I__1835 (
            .O(N__21806),
            .I(N__21803));
    Span4Mux_v I__1834 (
            .O(N__21803),
            .I(N__21800));
    Span4Mux_v I__1833 (
            .O(N__21800),
            .I(N__21797));
    Odrv4 I__1832 (
            .O(N__21797),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1831 (
            .O(N__21794),
            .I(N__21791));
    LocalMux I__1830 (
            .O(N__21791),
            .I(\pwm_generator_inst.un18_threshold_1_axb_0 ));
    InMux I__1829 (
            .O(N__21788),
            .I(N__21785));
    LocalMux I__1828 (
            .O(N__21785),
            .I(N__21782));
    Sp12to4 I__1827 (
            .O(N__21782),
            .I(N__21779));
    Span12Mux_s11_v I__1826 (
            .O(N__21779),
            .I(N__21776));
    Span12Mux_h I__1825 (
            .O(N__21776),
            .I(N__21773));
    Span12Mux_h I__1824 (
            .O(N__21773),
            .I(N__21770));
    Odrv12 I__1823 (
            .O(N__21770),
            .I(\pwm_generator_inst.O_0_1 ));
    InMux I__1822 (
            .O(N__21767),
            .I(N__21764));
    LocalMux I__1821 (
            .O(N__21764),
            .I(N__21761));
    Sp12to4 I__1820 (
            .O(N__21761),
            .I(N__21758));
    Span12Mux_s10_v I__1819 (
            .O(N__21758),
            .I(N__21755));
    Span12Mux_h I__1818 (
            .O(N__21755),
            .I(N__21752));
    Span12Mux_h I__1817 (
            .O(N__21752),
            .I(N__21749));
    Odrv12 I__1816 (
            .O(N__21749),
            .I(\pwm_generator_inst.O_0_0 ));
    InMux I__1815 (
            .O(N__21746),
            .I(N__21743));
    LocalMux I__1814 (
            .O(N__21743),
            .I(N__21740));
    Span4Mux_v I__1813 (
            .O(N__21740),
            .I(N__21737));
    Sp12to4 I__1812 (
            .O(N__21737),
            .I(N__21734));
    Span12Mux_h I__1811 (
            .O(N__21734),
            .I(N__21731));
    Span12Mux_h I__1810 (
            .O(N__21731),
            .I(N__21728));
    Span12Mux_v I__1809 (
            .O(N__21728),
            .I(N__21725));
    Odrv12 I__1808 (
            .O(N__21725),
            .I(\pwm_generator_inst.O_0_5 ));
    InMux I__1807 (
            .O(N__21722),
            .I(N__21719));
    LocalMux I__1806 (
            .O(N__21719),
            .I(N__21716));
    Sp12to4 I__1805 (
            .O(N__21716),
            .I(N__21713));
    Span12Mux_s5_v I__1804 (
            .O(N__21713),
            .I(N__21710));
    Span12Mux_h I__1803 (
            .O(N__21710),
            .I(N__21707));
    Span12Mux_h I__1802 (
            .O(N__21707),
            .I(N__21704));
    Odrv12 I__1801 (
            .O(N__21704),
            .I(\pwm_generator_inst.O_0_3 ));
    InMux I__1800 (
            .O(N__21701),
            .I(N__21698));
    LocalMux I__1799 (
            .O(N__21698),
            .I(N__21695));
    Span12Mux_s1_h I__1798 (
            .O(N__21695),
            .I(N__21692));
    Span12Mux_h I__1797 (
            .O(N__21692),
            .I(N__21689));
    Span12Mux_h I__1796 (
            .O(N__21689),
            .I(N__21686));
    Odrv12 I__1795 (
            .O(N__21686),
            .I(\pwm_generator_inst.O_0_4 ));
    InMux I__1794 (
            .O(N__21683),
            .I(N__21680));
    LocalMux I__1793 (
            .O(N__21680),
            .I(N__21677));
    Sp12to4 I__1792 (
            .O(N__21677),
            .I(N__21674));
    Span12Mux_v I__1791 (
            .O(N__21674),
            .I(N__21671));
    Span12Mux_h I__1790 (
            .O(N__21671),
            .I(N__21668));
    Span12Mux_h I__1789 (
            .O(N__21668),
            .I(N__21665));
    Odrv12 I__1788 (
            .O(N__21665),
            .I(\pwm_generator_inst.O_0_2 ));
    InMux I__1787 (
            .O(N__21662),
            .I(N__21659));
    LocalMux I__1786 (
            .O(N__21659),
            .I(N__21656));
    Span4Mux_v I__1785 (
            .O(N__21656),
            .I(N__21653));
    Sp12to4 I__1784 (
            .O(N__21653),
            .I(N__21650));
    Span12Mux_h I__1783 (
            .O(N__21650),
            .I(N__21647));
    Span12Mux_h I__1782 (
            .O(N__21647),
            .I(N__21644));
    Odrv12 I__1781 (
            .O(N__21644),
            .I(\pwm_generator_inst.O_0_6 ));
    IoInMux I__1780 (
            .O(N__21641),
            .I(N__21638));
    LocalMux I__1779 (
            .O(N__21638),
            .I(N__21635));
    IoSpan4Mux I__1778 (
            .O(N__21635),
            .I(N__21632));
    IoSpan4Mux I__1777 (
            .O(N__21632),
            .I(N__21629));
    Odrv4 I__1776 (
            .O(N__21629),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    IoInMux I__1775 (
            .O(N__21626),
            .I(N__21623));
    LocalMux I__1774 (
            .O(N__21623),
            .I(N__21620));
    Span4Mux_s3_v I__1773 (
            .O(N__21620),
            .I(N__21617));
    Span4Mux_h I__1772 (
            .O(N__21617),
            .I(N__21614));
    Sp12to4 I__1771 (
            .O(N__21614),
            .I(N__21611));
    Span12Mux_v I__1770 (
            .O(N__21611),
            .I(N__21608));
    Span12Mux_v I__1769 (
            .O(N__21608),
            .I(N__21605));
    Odrv12 I__1768 (
            .O(N__21605),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\pwm_generator_inst.un22_threshold_1_cry_7 ),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_18_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_23_0_));
    defparam IN_MUX_bfv_18_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_24_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_18_24_0_));
    defparam IN_MUX_bfv_18_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_25_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_18_25_0_));
    defparam IN_MUX_bfv_18_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_26_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_18_26_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\pwm_generator_inst.un5_threshold_add_1_cry_7 ),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(\pwm_generator_inst.un5_threshold_add_1_cry_15 ),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\pwm_generator_inst.un18_threshold_1_cry_7 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\pwm_generator_inst.un18_threshold_1_cry_15 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\pwm_generator_inst.un18_threshold_1_cry_23 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_3_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_12_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_30 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_7 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_15 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_23 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_30 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_10_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_2_0_));
    defparam IN_MUX_bfv_10_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_3_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_7 ),
            .carryinitout(bfn_10_3_0_));
    defparam IN_MUX_bfv_10_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_4_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_15 ),
            .carryinitout(bfn_10_4_0_));
    defparam IN_MUX_bfv_10_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_5_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_23 ),
            .carryinitout(bfn_10_5_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_30 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_7 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_15 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_8_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_23_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_23 ),
            .carryinitout(bfn_8_23_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_30 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_7 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_15 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_23 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_17_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_3_0_));
    defparam IN_MUX_bfv_17_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_4_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_4_0_));
    defparam IN_MUX_bfv_17_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_5_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_5_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_15 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_23 ),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_17_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_25_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_17_25_0_));
    defparam IN_MUX_bfv_17_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_26_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_17_26_0_));
    defparam IN_MUX_bfv_12_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_23_0_));
    defparam IN_MUX_bfv_12_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_24_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_12_24_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_15_24_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21626),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21641),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \phase_controller_inst1.stoper_tr.running_RNI6D081_0  (
            .USERSIGNALTOGLOBALBUFFER(N__29003),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst1.stoper_tr.un2_start_0_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.running_RNI96ON_0  (
            .USERSIGNALTOGLOBALBUFFER(N__24539),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un2_start_0_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__49010),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_163_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__42106),
            .CLKHFEN(N__42110),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__42218),
            .RGB2PWM(N__23027),
            .RGB1(rgb_g),
            .CURREN(N__42779),
            .RGB2(rgb_b),
            .RGB1PWM(N__23327),
            .RGB0PWM(N__53465),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__21794),
            .in2(_gnd_net_),
            .in3(N__21809),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__21938),
            .in2(_gnd_net_),
            .in3(N__21953),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_13_2  (
            .in0(N__21932),
            .in1(N__21917),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_13_3  (
            .in0(N__21911),
            .in1(N__21896),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__21875),
            .in2(_gnd_net_),
            .in3(N__21890),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__21854),
            .in2(_gnd_net_),
            .in3(N__21869),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__21833),
            .in2(_gnd_net_),
            .in3(N__21848),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__21815),
            .in2(_gnd_net_),
            .in3(N__21827),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__22085),
            .in2(_gnd_net_),
            .in3(N__22097),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__22064),
            .in2(_gnd_net_),
            .in3(N__22079),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__22043),
            .in2(_gnd_net_),
            .in3(N__22058),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_10 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__22022),
            .in2(_gnd_net_),
            .in3(N__22037),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__22001),
            .in2(_gnd_net_),
            .in3(N__22016),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_12 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__21980),
            .in2(_gnd_net_),
            .in3(N__21995),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_13 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__21959),
            .in2(_gnd_net_),
            .in3(N__21974),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_14 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__22172),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__22133),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__22223),
            .in2(_gnd_net_),
            .in3(N__22121),
            .lcout(\pwm_generator_inst.un22_threshold_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__22217),
            .in2(_gnd_net_),
            .in3(N__22118),
            .lcout(\pwm_generator_inst.un18_threshold1_18 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__23507),
            .in2(_gnd_net_),
            .in3(N__22115),
            .lcout(\pwm_generator_inst.un18_threshold1_19 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_18 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__22229),
            .in2(_gnd_net_),
            .in3(N__22112),
            .lcout(\pwm_generator_inst.un18_threshold1_20 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_19 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__22205),
            .in2(_gnd_net_),
            .in3(N__22109),
            .lcout(\pwm_generator_inst.un18_threshold1_21 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_20 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__22211),
            .in2(_gnd_net_),
            .in3(N__22106),
            .lcout(\pwm_generator_inst.un18_threshold1_22 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_21 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__23186),
            .in2(_gnd_net_),
            .in3(N__22103),
            .lcout(\pwm_generator_inst.un18_threshold1_23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_22 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__23141),
            .in2(_gnd_net_),
            .in3(N__22100),
            .lcout(\pwm_generator_inst.un18_threshold1_24 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__23333),
            .in2(_gnd_net_),
            .in3(N__22235),
            .lcout(\pwm_generator_inst.un18_threshold1_25 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_24 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_16_2 .LUT_INIT=16'b0110101010011010;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_16_2  (
            .in0(N__22556),
            .in1(N__23273),
            .in2(N__23899),
            .in3(N__22232),
            .lcout(\pwm_generator_inst.N_188_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_16_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23965),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23233),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_16_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23005),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23806),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23920),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_17_0 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__22199),
            .in2(N__22187),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_15 ),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_17_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__22163),
            .in2(N__22151),
            .in3(N__22124),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_16 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__22502),
            .in2(N__22490),
            .in3(N__22472),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__22469),
            .in2(N__22457),
            .in3(N__22436),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__22433),
            .in2(N__22421),
            .in3(N__22403),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__22400),
            .in2(N__22388),
            .in3(N__22370),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__22367),
            .in2(N__22352),
            .in3(N__22337),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__22334),
            .in2(N__22319),
            .in3(N__22304),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__22301),
            .in2(N__22286),
            .in3(N__22271),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0 ),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_18_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__22268),
            .in2(N__22253),
            .in3(N__22238),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_18_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__22604),
            .in2(N__22589),
            .in3(N__22574),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_18_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__23477),
            .in2(N__22571),
            .in3(N__22547),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_18_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__22544),
            .in2(N__23492),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_18_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__23481),
            .in2(N__22532),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_18_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__22517),
            .in2(N__23493),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_18_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__23485),
            .in2(N__23042),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_19_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__23357),
            .in2(_gnd_net_),
            .in3(N__22505),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_20_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(N__29879),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_20_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__22862),
            .in2(_gnd_net_),
            .in3(N__22829),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_20_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(N__41989),
            .in2(N__22826),
            .in3(N__22790),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_20_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_20_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_20_3  (
            .in0(_gnd_net_),
            .in1(N__22787),
            .in2(N__42095),
            .in3(N__22754),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_20_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(N__22751),
            .in2(_gnd_net_),
            .in3(N__22721),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_20_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_20_5  (
            .in0(_gnd_net_),
            .in1(N__22718),
            .in2(N__42096),
            .in3(N__22691),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_20_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_20_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_20_6  (
            .in0(_gnd_net_),
            .in1(N__22688),
            .in2(_gnd_net_),
            .in3(N__22655),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_20_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_20_7  (
            .in0(_gnd_net_),
            .in1(N__22652),
            .in2(_gnd_net_),
            .in3(N__22622),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_21_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_21_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36773),
            .in3(N__22607),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0 ),
            .ltout(),
            .carryin(bfn_1_21_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_21_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_21_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_21_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36722),
            .in3(N__22982),
            .lcout(\pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_21_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_21_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36665),
            .in3(N__22967),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_21_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_21_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_21_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36608),
            .in3(N__22952),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_21_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_21_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(N__37142),
            .in2(_gnd_net_),
            .in3(N__22937),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_21_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_21_5  (
            .in0(_gnd_net_),
            .in1(N__37106),
            .in2(_gnd_net_),
            .in3(N__22922),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_21_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_21_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_21_6  (
            .in0(_gnd_net_),
            .in1(N__37076),
            .in2(_gnd_net_),
            .in3(N__22907),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_21_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_21_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_21_7  (
            .in0(_gnd_net_),
            .in1(N__37037),
            .in2(_gnd_net_),
            .in3(N__22892),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_22_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(N__37001),
            .in2(_gnd_net_),
            .in3(N__22877),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7 ),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_22_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_22_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(N__36968),
            .in2(_gnd_net_),
            .in3(N__23078),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_22_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_22_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_22_2  (
            .in0(_gnd_net_),
            .in1(N__36932),
            .in2(_gnd_net_),
            .in3(N__23063),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_22_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(N__37334),
            .in2(_gnd_net_),
            .in3(N__23060),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_22_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_22_4  (
            .in0(N__37316),
            .in1(N__23057),
            .in2(N__36896),
            .in3(N__23045),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_22_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_22_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_22_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_22_7  (
            .in0(N__23494),
            .in1(N__23398),
            .in2(_gnd_net_),
            .in3(N__23380),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.N_112_i_i_LC_1_29_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_112_i_i_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_112_i_i_LC_1_29_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \phase_controller_inst1.N_112_i_i_LC_1_29_3  (
            .in0(N__26992),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53463),
            .lcout(N_112_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_2_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_2_13_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNITBL3_9_LC_2_13_1  (
            .in0(N__24048),
            .in1(N__24087),
            .in2(_gnd_net_),
            .in3(N__24222),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_2_13_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_2_13_4 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_2_LC_2_13_4  (
            .in0(N__23676),
            .in1(N__23631),
            .in2(N__23708),
            .in3(N__23135),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_2_13_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_2_13_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_6_LC_2_13_5  (
            .in0(N__23021),
            .in1(N__24126),
            .in2(N__23015),
            .in3(N__24184),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_13_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_13_6 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_13_6  (
            .in0(N__23108),
            .in1(N__23889),
            .in2(N__23129),
            .in3(N__23012),
            .lcout(\pwm_generator_inst.N_180_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_2_13_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_2_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIRPD2_0_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__23781),
            .in2(_gnd_net_),
            .in3(N__23754),
            .lcout(\pwm_generator_inst.un1_counterlto2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__23245),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__42190),
            .in2(N__23125),
            .in3(N__23099),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__23536),
            .in2(N__42342),
            .in3(N__23096),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__42194),
            .in2(N__23998),
            .in3(N__23093),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__23938),
            .in2(N__42343),
            .in3(N__23090),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__42198),
            .in2(N__23830),
            .in3(N__23087),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__23206),
            .in2(N__42344),
            .in3(N__23084),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__42202),
            .in2(N__23177),
            .in3(N__23081),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__23263),
            .in2(N__42189),
            .in3(N__23279),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23276),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_16_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_16_6  (
            .in0(N__23348),
            .in1(N__23885),
            .in2(N__23267),
            .in3(N__23252),
            .lcout(\pwm_generator_inst.N_187_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_16_7  (
            .in0(N__23884),
            .in1(N__23246),
            .in2(_gnd_net_),
            .in3(N__23234),
            .lcout(\pwm_generator_inst.N_179_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_17_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_17_0 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_17_0  (
            .in0(N__23195),
            .in1(N__23222),
            .in2(N__23213),
            .in3(N__23879),
            .lcout(\pwm_generator_inst.N_185_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_2_17_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_2_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23194),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_2_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_2_17_2 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_2_17_2  (
            .in0(N__23150),
            .in1(N__23176),
            .in2(N__23162),
            .in3(N__23880),
            .lcout(\pwm_generator_inst.N_186_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_2_17_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_2_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23149),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_2_17_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_2_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__23495),
            .in2(_gnd_net_),
            .in3(N__23432),
            .lcout(),
            .ltout(\pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_2_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_2_17_6 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_2_17_6  (
            .in0(N__23417),
            .in1(N__23405),
            .in2(N__23387),
            .in3(N__23384),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_2_17_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_2_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23344),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un8_start_stop_LC_2_30_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.un8_start_stop_LC_2_30_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un8_start_stop_LC_2_30_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.un8_start_stop_LC_2_30_0  (
            .in0(N__53464),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26996),
            .lcout(un8_start_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_3.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_2_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23318),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_3_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_3_12_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_3_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_3_12_0  (
            .in0(N__23588),
            .in1(N__23785),
            .in2(_gnd_net_),
            .in3(N__23291),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_3_12_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__53843),
            .ce(),
            .sr(N__53396));
    defparam \pwm_generator_inst.counter_1_LC_3_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_3_12_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_3_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_3_12_1  (
            .in0(N__23582),
            .in1(N__23758),
            .in2(_gnd_net_),
            .in3(N__23288),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__53843),
            .ce(),
            .sr(N__53396));
    defparam \pwm_generator_inst.counter_2_LC_3_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_3_12_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_3_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_3_12_2  (
            .in0(N__23589),
            .in1(N__23706),
            .in2(_gnd_net_),
            .in3(N__23285),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__53843),
            .ce(),
            .sr(N__53396));
    defparam \pwm_generator_inst.counter_3_LC_3_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_3_12_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_3_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_3_12_3  (
            .in0(N__23583),
            .in1(N__23677),
            .in2(_gnd_net_),
            .in3(N__23282),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__53843),
            .ce(),
            .sr(N__53396));
    defparam \pwm_generator_inst.counter_4_LC_3_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_3_12_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_3_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_3_12_4  (
            .in0(N__23590),
            .in1(N__23632),
            .in2(_gnd_net_),
            .in3(N__23606),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__53843),
            .ce(),
            .sr(N__53396));
    defparam \pwm_generator_inst.counter_5_LC_3_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_3_12_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_3_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_3_12_5  (
            .in0(N__23584),
            .in1(N__24223),
            .in2(_gnd_net_),
            .in3(N__23603),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__53843),
            .ce(),
            .sr(N__53396));
    defparam \pwm_generator_inst.counter_6_LC_3_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_3_12_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_3_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_3_12_6  (
            .in0(N__23591),
            .in1(N__24183),
            .in2(_gnd_net_),
            .in3(N__23600),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__53843),
            .ce(),
            .sr(N__53396));
    defparam \pwm_generator_inst.counter_7_LC_3_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_3_12_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_3_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_3_12_7  (
            .in0(N__23585),
            .in1(N__24127),
            .in2(_gnd_net_),
            .in3(N__23597),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__53843),
            .ce(),
            .sr(N__53396));
    defparam \pwm_generator_inst.counter_8_LC_3_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_3_13_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_3_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_3_13_0  (
            .in0(N__23587),
            .in1(N__24091),
            .in2(_gnd_net_),
            .in3(N__23594),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__53837),
            .ce(),
            .sr(N__53405));
    defparam \pwm_generator_inst.counter_9_LC_3_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_3_13_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_3_13_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_3_13_1  (
            .in0(N__24052),
            .in1(N__23586),
            .in2(_gnd_net_),
            .in3(N__23552),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53837),
            .ce(),
            .sr(N__53405));
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_3_14_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_3_14_0 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_3_14_0  (
            .in0(N__23549),
            .in1(N__23900),
            .in2(N__23525),
            .in3(N__23543),
            .lcout(\pwm_generator_inst.N_181_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_3_14_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_3_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23521),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_3_14_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_3_14_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_3_14_2  (
            .in0(N__24002),
            .in1(N__23981),
            .in2(N__23975),
            .in3(N__23902),
            .lcout(\pwm_generator_inst.N_182_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_3_14_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_3_14_4 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_3_14_4  (
            .in0(N__23954),
            .in1(N__23903),
            .in2(N__23948),
            .in3(N__23927),
            .lcout(\pwm_generator_inst.N_183_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_3_14_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_3_14_6 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_3_14_6  (
            .in0(N__23909),
            .in1(N__23901),
            .in2(N__23837),
            .in3(N__23813),
            .lcout(\pwm_generator_inst.N_184_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__23765),
            .in2(N__23795),
            .in3(N__23786),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_15_1  (
            .in0(N__23759),
            .in1(N__23723),
            .in2(N__23738),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__23684),
            .in2(N__23717),
            .in3(N__23707),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_15_3  (
            .in0(N__23678),
            .in1(N__23648),
            .in2(N__23657),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__23612),
            .in2(N__23642),
            .in3(N__23633),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_15_5  (
            .in0(N__24224),
            .in1(N__24191),
            .in2(N__24203),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_15_6  (
            .in0(N__24185),
            .in1(N__24149),
            .in2(N__24164),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__24107),
            .in2(N__24143),
            .in3(N__24128),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__24071),
            .in2(N__24101),
            .in3(N__24092),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__24032),
            .in2(N__24065),
            .in3(N__24053),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_3_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_3_16_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_3_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24026),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53817),
            .ce(),
            .sr(N__53415));
    defparam CONSTANT_ONE_LUT4_LC_3_21_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_3_21_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_3_21_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_3_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_4_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_4_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_15_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26351),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53824),
            .ce(N__24456),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_4_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_4_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_4_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_12_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26120),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53818),
            .ce(N__24448),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_5_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_14_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26372),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53819),
            .ce(N__24443),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_5_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_5_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_28_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27793),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53809),
            .ce(N__24447),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_5_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_5_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_2_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26045),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53801),
            .ce(N__24457),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_5_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_5_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_13_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26393),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53801),
            .ce(N__24457),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_17_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28499),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53794),
            .ce(N__24455),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__25866),
            .in2(_gnd_net_),
            .in3(N__24615),
            .lcout(\phase_controller_inst2.stoper_tr.un4_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_7_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_7_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_7_7_0 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_7_7_0  (
            .in0(N__26820),
            .in1(N__24569),
            .in2(N__26797),
            .in3(N__24620),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53847),
            .ce(),
            .sr(N__53344));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_7_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_7_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_7_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_7_7_1  (
            .in0(N__24621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53847),
            .ce(),
            .sr(N__53344));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_8_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_7_8_1  (
            .in0(N__41094),
            .in1(N__41133),
            .in2(_gnd_net_),
            .in3(N__38558),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53844),
            .ce(),
            .sr(N__53348));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_7_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_7_9_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_7_9_2  (
            .in0(N__25874),
            .in1(N__53460),
            .in2(_gnd_net_),
            .in3(N__24623),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_7_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_7_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25875),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_7_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_7_10_2 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_7_10_2 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.state_4_LC_7_10_2  (
            .in0(N__26884),
            .in1(N__26910),
            .in2(_gnd_net_),
            .in3(N__26976),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53830),
            .ce(),
            .sr(N__53363));
    defparam \phase_controller_inst1.start_flag_LC_7_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_flag_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_flag_LC_7_10_3 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \phase_controller_inst1.start_flag_LC_7_10_3  (
            .in0(N__26975),
            .in1(_gnd_net_),
            .in2(N__26917),
            .in3(N__26883),
            .lcout(\phase_controller_inst1.start_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53830),
            .ce(),
            .sr(N__53363));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_11_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_11_0  (
            .in0(N__24511),
            .in1(N__24961),
            .in2(N__24322),
            .in3(N__24706),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_11_2 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_11_2  (
            .in0(N__24512),
            .in1(N__24960),
            .in2(N__24323),
            .in3(N__24705),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_11_4 .LUT_INIT=16'b0010001010110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_11_4  (
            .in0(N__24233),
            .in1(N__24924),
            .in2(N__24484),
            .in3(N__24943),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_11_6 .LUT_INIT=16'b1011001010111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_11_6  (
            .in0(N__24232),
            .in1(N__24925),
            .in2(N__24485),
            .in3(N__24942),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30191),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53825),
            .ce(N__24406),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_7_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_7_12_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_7_12_0  (
            .in0(N__24524),
            .in1(N__24889),
            .in2(N__24269),
            .in3(N__24907),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_7_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_7_12_2 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_7_12_2  (
            .in0(N__24523),
            .in1(N__24888),
            .in2(N__24268),
            .in3(N__24906),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_7_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_7_12_4 .LUT_INIT=16'b0000101010001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_7_12_4  (
            .in0(N__24335),
            .in1(N__24497),
            .in2(N__24854),
            .in3(N__24871),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_7_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_7_12_6 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_7_12_6  (
            .in0(N__24334),
            .in1(N__24496),
            .in2(N__24853),
            .in3(N__24870),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_13_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_13_0  (
            .in0(N__33116),
            .in1(N__41053),
            .in2(_gnd_net_),
            .in3(N__31772),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(elapsed_time_ns_1_RNI0CQBB_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_13_1 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_13_1  (
            .in0(N__41020),
            .in1(_gnd_net_),
            .in2(N__24245),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53810),
            .ce(N__24407),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_13_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_13_2  (
            .in0(N__32777),
            .in1(N__24242),
            .in2(_gnd_net_),
            .in3(N__31773),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(elapsed_time_ns_1_RNI1BOBB_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_7_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_7_13_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24236),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_13_4  (
            .in0(N__26089),
            .in1(N__32963),
            .in2(_gnd_net_),
            .in3(N__31774),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_7_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_7_14_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_7_14_0  (
            .in0(N__24287),
            .in1(N__24785),
            .in2(N__24815),
            .in3(N__24278),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_7_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_7_14_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_7_14_2  (
            .in0(N__24286),
            .in1(N__24784),
            .in2(N__24814),
            .in3(N__24277),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_14_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_14_4  (
            .in0(N__24296),
            .in1(N__24731),
            .in2(N__24761),
            .in3(N__24305),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_7_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_7_14_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_7_14_6  (
            .in0(N__24295),
            .in1(N__24730),
            .in2(N__24760),
            .in3(N__24304),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_7_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_7_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_19_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26267),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53802),
            .ce(N__24437),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26060),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53795),
            .ce(N__24439),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26138),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53795),
            .ce(N__24439),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_15_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_15_2  (
            .in0(N__26203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53795),
            .ce(N__24439),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_7_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_7_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_18_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26288),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53795),
            .ce(N__24439),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_7_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_7_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_16_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26330),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53795),
            .ce(N__24439),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_7_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_7_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_17_LC_7_15_5  (
            .in0(N__26309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53795),
            .ce(N__24439),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_7_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_7_15_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_27_LC_7_15_6  (
            .in0(N__26420),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53795),
            .ce(N__24439),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26027),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53795),
            .ce(N__24439),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26008),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53788),
            .ce(N__24438),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26236),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53788),
            .ce(N__24438),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26218),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53788),
            .ce(N__24438),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30224),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53788),
            .ce(N__24438),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26186),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53788),
            .ce(N__24438),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26153),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53788),
            .ce(N__24438),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_7_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_7_17_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__26059),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53786),
            .ce(N__40956),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_7_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_7_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_11_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26134),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53786),
            .ce(N__40956),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_7_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_7_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_12_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26113),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53786),
            .ce(N__40956),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_7_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_7_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_13_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26386),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53786),
            .ce(N__40956),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_7_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_7_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_14_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26365),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53786),
            .ce(N__40956),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_7_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_7_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_15_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26344),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53786),
            .ce(N__40956),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_7_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_7_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_2_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26041),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53786),
            .ce(N__40956),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_7_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_7_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_3_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26026),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53786),
            .ce(N__40956),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_7_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_7_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_4_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26012),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53783),
            .ce(N__40955),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_7_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_7_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_5_LC_7_18_1  (
            .in0(N__26240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53783),
            .ce(N__40955),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_7_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_7_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_6_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26222),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53783),
            .ce(N__40955),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_7_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_7_18_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_7_LC_7_18_3  (
            .in0(N__26204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53783),
            .ce(N__40955),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_7_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_7_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_8_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26185),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53783),
            .ce(N__40955),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_7_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_7_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_9_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26167),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53783),
            .ce(N__40955),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_7_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_7_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_10_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26152),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53783),
            .ce(N__40955),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_7_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_7_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_24_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28510),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53782),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30238),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53782),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_7_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_7_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_26_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28465),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53782),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26171),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53782),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30205),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53782),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_7_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_7_20_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_7_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_16_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26329),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53778),
            .ce(N__40954),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_7_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_7_20_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_7_20_2  (
            .in0(N__28651),
            .in1(N__28640),
            .in2(N__28619),
            .in3(N__28585),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_7_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_7_20_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_7_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_17_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26308),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53778),
            .ce(N__40954),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_20_4 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_7_20_4  (
            .in0(N__26483),
            .in1(N__24557),
            .in2(N__26510),
            .in3(N__24548),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_7_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_7_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_18_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26284),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53778),
            .ce(N__40954),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_7_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_7_20_6 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_7_20_6  (
            .in0(N__26482),
            .in1(N__24556),
            .in2(N__26509),
            .in3(N__24547),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_7_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_7_20_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_7_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_19_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26263),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53778),
            .ce(N__40954),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_7_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_7_22_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_7_22_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_27_LC_7_22_6  (
            .in0(N__26416),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53766),
            .ce(N__40937),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_5_2 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_8_5_2  (
            .in0(N__24582),
            .in1(N__24622),
            .in2(_gnd_net_),
            .in3(N__25873),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_8_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_8_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_8_6_0 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst2.state_0_LC_8_6_0  (
            .in0(N__26576),
            .in1(N__26787),
            .in2(N__26600),
            .in3(N__26834),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53848),
            .ce(),
            .sr(N__53339));
    defparam \phase_controller_inst2.state_3_LC_8_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_8_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_8_6_1 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \phase_controller_inst2.state_3_LC_8_6_1  (
            .in0(N__24652),
            .in1(N__26970),
            .in2(N__24640),
            .in3(N__26564),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53848),
            .ce(),
            .sr(N__53339));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_8_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_8_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_8_6_3 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_8_6_3  (
            .in0(N__26595),
            .in1(N__24583),
            .in2(N__24662),
            .in3(N__25828),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53848),
            .ce(),
            .sr(N__53339));
    defparam \phase_controller_inst2.state_4_LC_8_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_4_LC_8_6_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst2.state_4_LC_8_6_5 .LUT_INIT=16'b1010000010101010;
    LogicCell40 \phase_controller_inst2.state_4_LC_8_6_5  (
            .in0(N__24653),
            .in1(_gnd_net_),
            .in2(N__24641),
            .in3(N__26971),
            .lcout(\phase_controller_inst2.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53848),
            .ce(),
            .sr(N__53339));
    defparam \phase_controller_inst2.start_flag_LC_8_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_flag_LC_8_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_flag_LC_8_6_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \phase_controller_inst2.start_flag_LC_8_6_6  (
            .in0(N__26969),
            .in1(N__24651),
            .in2(_gnd_net_),
            .in3(N__24639),
            .lcout(\phase_controller_inst2.start_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53848),
            .ce(),
            .sr(N__53339));
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_8_6_7 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_8_6_7  (
            .in0(N__24619),
            .in1(N__24584),
            .in2(N__25876),
            .in3(N__25829),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53848),
            .ce(),
            .sr(N__53339));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__26723),
            .in2(_gnd_net_),
            .in3(N__26651),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_8_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_8_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__26698),
            .in2(_gnd_net_),
            .in3(N__30675),
            .lcout(\phase_controller_inst2.stoper_hc.un4_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_8_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_8_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_0_LC_8_8_0  (
            .in0(N__25259),
            .in1(N__25135),
            .in2(N__25808),
            .in3(N__25807),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_0 ),
            .clk(N__53838),
            .ce(N__25157),
            .sr(N__53345));
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_8_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_8_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_8_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_1_LC_8_8_1  (
            .in0(N__25267),
            .in1(N__25102),
            .in2(_gnd_net_),
            .in3(N__24563),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_1 ),
            .clk(N__53838),
            .ce(N__25157),
            .sr(N__53345));
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_8_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_8_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_2_LC_8_8_2  (
            .in0(N__25260),
            .in1(N__25066),
            .in2(_gnd_net_),
            .in3(N__24560),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_2 ),
            .clk(N__53838),
            .ce(N__25157),
            .sr(N__53345));
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_8_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_8_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_8_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_3_LC_8_8_3  (
            .in0(N__25268),
            .in1(N__25027),
            .in2(_gnd_net_),
            .in3(N__24689),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_3 ),
            .clk(N__53838),
            .ce(N__25157),
            .sr(N__53345));
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_8_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_8_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_8_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_4_LC_8_8_4  (
            .in0(N__25261),
            .in1(N__24988),
            .in2(_gnd_net_),
            .in3(N__24686),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_4 ),
            .clk(N__53838),
            .ce(N__25157),
            .sr(N__53345));
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_8_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_8_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_5_LC_8_8_5  (
            .in0(N__25269),
            .in1(N__25546),
            .in2(_gnd_net_),
            .in3(N__24683),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_5 ),
            .clk(N__53838),
            .ce(N__25157),
            .sr(N__53345));
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_8_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_8_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_6_LC_8_8_6  (
            .in0(N__25262),
            .in1(N__25495),
            .in2(_gnd_net_),
            .in3(N__24680),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_6 ),
            .clk(N__53838),
            .ce(N__25157),
            .sr(N__53345));
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_8_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_8_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_8_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_7_LC_8_8_7  (
            .in0(N__25270),
            .in1(N__25456),
            .in2(_gnd_net_),
            .in3(N__24677),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_7 ),
            .clk(N__53838),
            .ce(N__25157),
            .sr(N__53345));
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_8_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_8_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_8_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_8_LC_8_9_0  (
            .in0(N__25258),
            .in1(N__25432),
            .in2(_gnd_net_),
            .in3(N__24674),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_8 ),
            .clk(N__53831),
            .ce(N__25158),
            .sr(N__53349));
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_8_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_8_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_9_LC_8_9_1  (
            .in0(N__25274),
            .in1(N__25384),
            .in2(_gnd_net_),
            .in3(N__24671),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_9 ),
            .clk(N__53831),
            .ce(N__25158),
            .sr(N__53349));
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_8_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_8_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_10_LC_8_9_2  (
            .in0(N__25255),
            .in1(N__25348),
            .in2(_gnd_net_),
            .in3(N__24668),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_10 ),
            .clk(N__53831),
            .ce(N__25158),
            .sr(N__53349));
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_8_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_8_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_11_LC_8_9_3  (
            .in0(N__25271),
            .in1(N__25312),
            .in2(_gnd_net_),
            .in3(N__24665),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_11 ),
            .clk(N__53831),
            .ce(N__25158),
            .sr(N__53349));
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_8_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_8_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_12_LC_8_9_4  (
            .in0(N__25256),
            .in1(N__25771),
            .in2(_gnd_net_),
            .in3(N__24827),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_12 ),
            .clk(N__53831),
            .ce(N__25158),
            .sr(N__53349));
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_8_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_8_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_13_LC_8_9_5  (
            .in0(N__25272),
            .in1(N__25747),
            .in2(_gnd_net_),
            .in3(N__24824),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_13 ),
            .clk(N__53831),
            .ce(N__25158),
            .sr(N__53349));
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_8_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_8_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_14_LC_8_9_6  (
            .in0(N__25257),
            .in1(N__25708),
            .in2(_gnd_net_),
            .in3(N__24821),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_14 ),
            .clk(N__53831),
            .ce(N__25158),
            .sr(N__53349));
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_8_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_8_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_15_LC_8_9_7  (
            .in0(N__25273),
            .in1(N__25669),
            .in2(_gnd_net_),
            .in3(N__24818),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_15 ),
            .clk(N__53831),
            .ce(N__25158),
            .sr(N__53349));
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_8_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_8_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_16_LC_8_10_0  (
            .in0(N__25283),
            .in1(N__24802),
            .in2(_gnd_net_),
            .in3(N__24788),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_16 ),
            .clk(N__53826),
            .ce(N__25159),
            .sr(N__53357));
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_8_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_8_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_17_LC_8_10_1  (
            .in0(N__25263),
            .in1(N__24778),
            .in2(_gnd_net_),
            .in3(N__24764),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_17 ),
            .clk(N__53826),
            .ce(N__25159),
            .sr(N__53357));
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_8_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_8_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_18_LC_8_10_2  (
            .in0(N__25284),
            .in1(N__24748),
            .in2(_gnd_net_),
            .in3(N__24734),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_18 ),
            .clk(N__53826),
            .ce(N__25159),
            .sr(N__53357));
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_8_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_8_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_19_LC_8_10_3  (
            .in0(N__25264),
            .in1(N__24724),
            .in2(_gnd_net_),
            .in3(N__24710),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_19 ),
            .clk(N__53826),
            .ce(N__25159),
            .sr(N__53357));
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_8_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_8_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_20_LC_8_10_4  (
            .in0(N__25285),
            .in1(N__24707),
            .in2(_gnd_net_),
            .in3(N__24692),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_20 ),
            .clk(N__53826),
            .ce(N__25159),
            .sr(N__53357));
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_8_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_8_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_21_LC_8_10_5  (
            .in0(N__25265),
            .in1(N__24962),
            .in2(_gnd_net_),
            .in3(N__24947),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_21 ),
            .clk(N__53826),
            .ce(N__25159),
            .sr(N__53357));
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_8_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_8_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_22_LC_8_10_6  (
            .in0(N__25286),
            .in1(N__24944),
            .in2(_gnd_net_),
            .in3(N__24929),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_22 ),
            .clk(N__53826),
            .ce(N__25159),
            .sr(N__53357));
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_8_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_8_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_23_LC_8_10_7  (
            .in0(N__25266),
            .in1(N__24926),
            .in2(_gnd_net_),
            .in3(N__24911),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_23 ),
            .clk(N__53826),
            .ce(N__25159),
            .sr(N__53357));
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_8_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_8_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_24_LC_8_11_0  (
            .in0(N__25275),
            .in1(N__24908),
            .in2(_gnd_net_),
            .in3(N__24893),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_24 ),
            .clk(N__53820),
            .ce(N__25160),
            .sr(N__53364));
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_8_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_8_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_25_LC_8_11_1  (
            .in0(N__25279),
            .in1(N__24890),
            .in2(_gnd_net_),
            .in3(N__24875),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_25 ),
            .clk(N__53820),
            .ce(N__25160),
            .sr(N__53364));
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_8_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_8_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_26_LC_8_11_2  (
            .in0(N__25276),
            .in1(N__24872),
            .in2(_gnd_net_),
            .in3(N__24857),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_26 ),
            .clk(N__53820),
            .ce(N__25160),
            .sr(N__53364));
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_8_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_8_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_27_LC_8_11_3  (
            .in0(N__25280),
            .in1(N__24852),
            .in2(_gnd_net_),
            .in3(N__24833),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_27 ),
            .clk(N__53820),
            .ce(N__25160),
            .sr(N__53364));
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_8_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_8_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_28_LC_8_11_4  (
            .in0(N__25277),
            .in1(N__25900),
            .in2(_gnd_net_),
            .in3(N__24830),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_28 ),
            .clk(N__53820),
            .ce(N__25160),
            .sr(N__53364));
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_8_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_8_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_29_LC_8_11_5  (
            .in0(N__25281),
            .in1(N__25924),
            .in2(_gnd_net_),
            .in3(N__25292),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_29 ),
            .clk(N__53820),
            .ce(N__25160),
            .sr(N__53364));
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_8_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_8_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_30_LC_8_11_6  (
            .in0(N__25278),
            .in1(N__34086),
            .in2(_gnd_net_),
            .in3(N__25289),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_29 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_30 ),
            .clk(N__53820),
            .ce(N__25160),
            .sr(N__53364));
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_8_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_8_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_31_LC_8_11_7  (
            .in0(N__25282),
            .in1(N__34116),
            .in2(_gnd_net_),
            .in3(N__25163),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53820),
            .ce(N__25160),
            .sr(N__53364));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_8_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_8_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__25142),
            .in2(N__25121),
            .in3(N__25136),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_0 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_8_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_8_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__25112),
            .in2(N__25088),
            .in3(N__25103),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_8_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_8_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__25079),
            .in2(N__25052),
            .in3(N__25067),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_8_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_8_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__25040),
            .in2(N__25013),
            .in3(N__25028),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_8_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_8_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__25004),
            .in2(N__24974),
            .in3(N__24992),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_8_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_8_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_8_12_5  (
            .in0(N__25547),
            .in1(N__25532),
            .in2(N__25520),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_8_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_8_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__25511),
            .in2(N__25481),
            .in3(N__25499),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_8_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_8_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__25469),
            .in2(N__25442),
            .in3(N__25460),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_8_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_8_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_8_13_0  (
            .in0(N__25433),
            .in1(N__25418),
            .in2(N__25406),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_8 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_8_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_8_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__25397),
            .in2(N__25370),
            .in3(N__25385),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_8_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_8_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__25361),
            .in2(N__25334),
            .in3(N__25349),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_8_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_8_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__25298),
            .in2(N__25325),
            .in3(N__25313),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_8_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_8_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__25784),
            .in2(N__25757),
            .in3(N__25772),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_8_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_8_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_8_13_5  (
            .in0(N__25748),
            .in1(N__25733),
            .in2(N__25721),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_8_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_8_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_8_13_6  (
            .in0(N__25709),
            .in1(N__25694),
            .in2(N__25682),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_8_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_8_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_8_13_7  (
            .in0(N__25673),
            .in1(N__25640),
            .in2(N__25655),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_8_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_8_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__25634),
            .in2(N__25628),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_8_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_8_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(N__25616),
            .in2(N__25610),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_8_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_8_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__25598),
            .in2(N__25586),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_8_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_8_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__25571),
            .in2(N__25562),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_8_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_8_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__25994),
            .in2(N__25985),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_8_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_8_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__25970),
            .in2(N__25961),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_8_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_8_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__25886),
            .in2(N__25943),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_8_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_8_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__34043),
            .in2(N__26075),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_8_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_8_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25946),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_8_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_8_15_1 .LUT_INIT=16'b0101111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_8_15_1  (
            .in0(N__25931),
            .in1(_gnd_net_),
            .in2(N__25910),
            .in3(N__34062),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_8_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_8_15_2 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_8_15_2  (
            .in0(N__34061),
            .in1(N__25930),
            .in2(_gnd_net_),
            .in3(N__25906),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_8_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_8_15_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__25880),
            .in2(_gnd_net_),
            .in3(N__25819),
            .lcout(\phase_controller_inst2.stoper_tr.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_8_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_8_15_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_8_15_4  (
            .in0(N__26099),
            .in1(N__32753),
            .in2(_gnd_net_),
            .in3(N__31787),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(elapsed_time_ns_1_RNI2COBB_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_15_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26093),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_8_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_8_15_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__26090),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_8_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_8_15_7 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_8_15_7  (
            .in0(N__34124),
            .in1(N__34097),
            .in2(_gnd_net_),
            .in3(N__34063),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__26066),
            .in2(N__41016),
            .in3(N__41073),
            .lcout(\phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_16_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_16_1  (
            .in0(N__27245),
            .in1(N__27241),
            .in2(N__42595),
            .in3(N__26048),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_1),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_16_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_16_2  (
            .in0(N__27221),
            .in1(N__27220),
            .in2(N__42599),
            .in3(N__26030),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_2),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_16_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_16_3  (
            .in0(N__27199),
            .in1(N__27200),
            .in2(N__42596),
            .in3(N__26015),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_3),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_16_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_16_4  (
            .in0(N__27170),
            .in1(N__27166),
            .in2(N__42600),
            .in3(N__25997),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_4),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_16_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_16_5  (
            .in0(N__27145),
            .in1(N__27146),
            .in2(N__42597),
            .in3(N__26225),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_5),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_16_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_16_6  (
            .in0(N__27125),
            .in1(N__27124),
            .in2(N__42601),
            .in3(N__26207),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_6),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_16_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_16_7  (
            .in0(N__27110),
            .in1(N__27109),
            .in2(N__42598),
            .in3(N__26189),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_7),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_17_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_17_0  (
            .in0(N__27095),
            .in1(N__27094),
            .in2(N__42362),
            .in3(N__26174),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_8),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_17_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_17_1  (
            .in0(N__27434),
            .in1(N__27430),
            .in2(N__42359),
            .in3(N__26156),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_9),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_17_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_17_2  (
            .in0(N__27410),
            .in1(N__27406),
            .in2(N__42363),
            .in3(N__26141),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_10),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_17_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_17_3  (
            .in0(N__27373),
            .in1(N__27374),
            .in2(N__42356),
            .in3(N__26123),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_11),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_17_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_17_4  (
            .in0(N__27344),
            .in1(N__27340),
            .in2(N__42360),
            .in3(N__26102),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_12),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_17_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_17_5  (
            .in0(N__27319),
            .in1(N__27320),
            .in2(N__42357),
            .in3(N__26375),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_13),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_17_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_17_6  (
            .in0(N__27299),
            .in1(N__27298),
            .in2(N__42361),
            .in3(N__26354),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_14),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_17_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_17_7  (
            .in0(N__27284),
            .in1(N__27283),
            .in2(N__42358),
            .in3(N__26333),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_15),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_18_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_18_0  (
            .in0(N__27268),
            .in1(N__27269),
            .in2(N__42452),
            .in3(N__26312),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_16),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_18_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_18_1  (
            .in0(N__27632),
            .in1(N__27628),
            .in2(N__42223),
            .in3(N__26291),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_17),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_18_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_18_2  (
            .in0(N__27599),
            .in1(N__27595),
            .in2(N__42453),
            .in3(N__26270),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_18),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_18_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_18_3  (
            .in0(N__27574),
            .in1(N__27575),
            .in2(N__42224),
            .in3(N__26249),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_19),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_18_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_18_4  (
            .in0(N__27548),
            .in1(N__27544),
            .in2(N__42454),
            .in3(N__26246),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_20),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_18_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_18_5  (
            .in0(N__27526),
            .in1(N__27527),
            .in2(N__42225),
            .in3(N__26243),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_21),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_18_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_18_6  (
            .in0(N__27506),
            .in1(N__27505),
            .in2(N__42455),
            .in3(N__26435),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_22),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_18_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_18_7  (
            .in0(N__27491),
            .in1(N__27490),
            .in2(N__42226),
            .in3(N__26432),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_23),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_19_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_19_0  (
            .in0(N__27476),
            .in1(N__27475),
            .in2(N__42219),
            .in3(N__26429),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_24),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_19_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_19_1  (
            .in0(N__27455),
            .in1(N__27451),
            .in2(N__42221),
            .in3(N__26426),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_25),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_19_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_19_2  (
            .in0(N__27851),
            .in1(N__27847),
            .in2(N__42220),
            .in3(N__26423),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_26),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_19_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_19_3  (
            .in0(N__27826),
            .in1(N__27827),
            .in2(N__42222),
            .in3(N__26402),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_27),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26399),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_8_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_8_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_0_LC_8_20_0  (
            .in0(N__28827),
            .in1(N__27757),
            .in2(N__28352),
            .in3(N__28351),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_0 ),
            .clk(N__53774),
            .ce(N__26627),
            .sr(N__53413));
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_8_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_8_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_8_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_1_LC_8_20_1  (
            .in0(N__28831),
            .in1(N__27721),
            .in2(_gnd_net_),
            .in3(N__26396),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_1 ),
            .clk(N__53774),
            .ce(N__26627),
            .sr(N__53413));
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_8_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_8_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_8_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_2_LC_8_20_2  (
            .in0(N__28828),
            .in1(N__27682),
            .in2(_gnd_net_),
            .in3(N__26462),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_2 ),
            .clk(N__53774),
            .ce(N__26627),
            .sr(N__53413));
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_8_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_8_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_3_LC_8_20_3  (
            .in0(N__28832),
            .in1(N__27646),
            .in2(_gnd_net_),
            .in3(N__26459),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_3 ),
            .clk(N__53774),
            .ce(N__26627),
            .sr(N__53413));
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_8_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_8_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_8_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_4_LC_8_20_4  (
            .in0(N__28829),
            .in1(N__28093),
            .in2(_gnd_net_),
            .in3(N__26456),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_4 ),
            .clk(N__53774),
            .ce(N__26627),
            .sr(N__53413));
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_8_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_8_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_8_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_5_LC_8_20_5  (
            .in0(N__28833),
            .in1(N__28066),
            .in2(_gnd_net_),
            .in3(N__26453),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_5 ),
            .clk(N__53774),
            .ce(N__26627),
            .sr(N__53413));
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_8_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_8_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_8_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_6_LC_8_20_6  (
            .in0(N__28830),
            .in1(N__28033),
            .in2(_gnd_net_),
            .in3(N__26450),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_6 ),
            .clk(N__53774),
            .ce(N__26627),
            .sr(N__53413));
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_8_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_8_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_8_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_7_LC_8_20_7  (
            .in0(N__28834),
            .in1(N__27997),
            .in2(_gnd_net_),
            .in3(N__26447),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_7 ),
            .clk(N__53774),
            .ce(N__26627),
            .sr(N__53413));
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_8_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_8_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_8_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_8_LC_8_21_0  (
            .in0(N__28813),
            .in1(N__27946),
            .in2(_gnd_net_),
            .in3(N__26444),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_8 ),
            .clk(N__53767),
            .ce(N__26626),
            .sr(N__53416));
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_8_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_8_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_9_LC_8_21_1  (
            .in0(N__28838),
            .in1(N__27913),
            .in2(_gnd_net_),
            .in3(N__26441),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_9 ),
            .clk(N__53767),
            .ce(N__26626),
            .sr(N__53416));
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_8_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_8_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_10_LC_8_21_2  (
            .in0(N__28810),
            .in1(N__27874),
            .in2(_gnd_net_),
            .in3(N__26438),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_10 ),
            .clk(N__53767),
            .ce(N__26626),
            .sr(N__53416));
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_8_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_8_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_11_LC_8_21_3  (
            .in0(N__28835),
            .in1(N__28315),
            .in2(_gnd_net_),
            .in3(N__26531),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_11 ),
            .clk(N__53767),
            .ce(N__26626),
            .sr(N__53416));
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_8_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_8_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_8_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_12_LC_8_21_4  (
            .in0(N__28811),
            .in1(N__28276),
            .in2(_gnd_net_),
            .in3(N__26528),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_12 ),
            .clk(N__53767),
            .ce(N__26626),
            .sr(N__53416));
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_8_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_8_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_8_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_13_LC_8_21_5  (
            .in0(N__28836),
            .in1(N__28255),
            .in2(_gnd_net_),
            .in3(N__26525),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_13 ),
            .clk(N__53767),
            .ce(N__26626),
            .sr(N__53416));
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_8_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_8_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_8_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_14_LC_8_21_6  (
            .in0(N__28812),
            .in1(N__28219),
            .in2(_gnd_net_),
            .in3(N__26522),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_14 ),
            .clk(N__53767),
            .ce(N__26626),
            .sr(N__53416));
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_8_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_8_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_8_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_15_LC_8_21_7  (
            .in0(N__28837),
            .in1(N__28183),
            .in2(_gnd_net_),
            .in3(N__26519),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_15 ),
            .clk(N__53767),
            .ce(N__26626),
            .sr(N__53416));
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_8_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_8_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_8_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_16_LC_8_22_0  (
            .in0(N__28806),
            .in1(N__28614),
            .in2(_gnd_net_),
            .in3(N__26516),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_16 ),
            .clk(N__53763),
            .ce(N__26625),
            .sr(N__53417));
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_8_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_8_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_8_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_17_LC_8_22_1  (
            .in0(N__28814),
            .in1(N__28639),
            .in2(_gnd_net_),
            .in3(N__26513),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_17 ),
            .clk(N__53763),
            .ce(N__26625),
            .sr(N__53417));
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_8_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_8_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_8_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_18_LC_8_22_2  (
            .in0(N__28807),
            .in1(N__26502),
            .in2(_gnd_net_),
            .in3(N__26486),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_18 ),
            .clk(N__53763),
            .ce(N__26625),
            .sr(N__53417));
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_8_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_8_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_8_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_19_LC_8_22_3  (
            .in0(N__28815),
            .in1(N__26481),
            .in2(_gnd_net_),
            .in3(N__26465),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_19 ),
            .clk(N__53763),
            .ce(N__26625),
            .sr(N__53417));
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_8_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_8_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_8_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_20_LC_8_22_4  (
            .in0(N__28808),
            .in1(N__30432),
            .in2(_gnd_net_),
            .in3(N__26558),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_20 ),
            .clk(N__53763),
            .ce(N__26625),
            .sr(N__53417));
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_8_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_8_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_8_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_21_LC_8_22_5  (
            .in0(N__28816),
            .in1(N__30480),
            .in2(_gnd_net_),
            .in3(N__26555),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_21 ),
            .clk(N__53763),
            .ce(N__26625),
            .sr(N__53417));
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_8_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_8_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_8_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_22_LC_8_22_6  (
            .in0(N__28809),
            .in1(N__30339),
            .in2(_gnd_net_),
            .in3(N__26552),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_22 ),
            .clk(N__53763),
            .ce(N__26625),
            .sr(N__53417));
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_8_22_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_8_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_8_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_23_LC_8_22_7  (
            .in0(N__28817),
            .in1(N__30367),
            .in2(_gnd_net_),
            .in3(N__26549),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_23 ),
            .clk(N__53763),
            .ce(N__26625),
            .sr(N__53417));
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_8_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_8_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_8_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_24_LC_8_23_0  (
            .in0(N__28780),
            .in1(N__28879),
            .in2(_gnd_net_),
            .in3(N__26546),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_23_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_24 ),
            .clk(N__53756),
            .ce(N__26624),
            .sr(N__53418));
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_8_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_8_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_8_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_25_LC_8_23_1  (
            .in0(N__28784),
            .in1(N__28912),
            .in2(_gnd_net_),
            .in3(N__26543),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_25 ),
            .clk(N__53756),
            .ce(N__26624),
            .sr(N__53418));
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_8_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_8_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_8_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_26_LC_8_23_2  (
            .in0(N__28781),
            .in1(N__28409),
            .in2(_gnd_net_),
            .in3(N__26540),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_26 ),
            .clk(N__53756),
            .ce(N__26624),
            .sr(N__53418));
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_8_23_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_8_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_8_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_27_LC_8_23_3  (
            .in0(N__28785),
            .in1(N__28451),
            .in2(_gnd_net_),
            .in3(N__26537),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_27 ),
            .clk(N__53756),
            .ce(N__26624),
            .sr(N__53418));
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_8_23_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_8_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_8_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_28_LC_8_23_4  (
            .in0(N__28782),
            .in1(N__28561),
            .in2(_gnd_net_),
            .in3(N__26534),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_28 ),
            .clk(N__53756),
            .ce(N__26624),
            .sr(N__53418));
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_8_23_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_8_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_8_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_29_LC_8_23_5  (
            .in0(N__28786),
            .in1(N__28545),
            .in2(_gnd_net_),
            .in3(N__26636),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_29 ),
            .clk(N__53756),
            .ce(N__26624),
            .sr(N__53418));
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_8_23_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_8_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_8_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_30_LC_8_23_6  (
            .in0(N__28783),
            .in1(N__28988),
            .in2(_gnd_net_),
            .in3(N__26633),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_30 ),
            .clk(N__53756),
            .ce(N__26624),
            .sr(N__53418));
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_8_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_8_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_8_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_31_LC_8_23_7  (
            .in0(N__28787),
            .in1(N__28943),
            .in2(_gnd_net_),
            .in3(N__26630),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53756),
            .ce(N__26624),
            .sr(N__53418));
    defparam \phase_controller_inst2.S2_LC_8_27_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_27_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_8_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26798),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53735),
            .ce(),
            .sr(N__53423));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_9_3_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_9_3_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_9_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30684),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_5_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_5_1  (
            .in0(N__30683),
            .in1(N__26678),
            .in2(_gnd_net_),
            .in3(N__26707),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_6  (
            .in0(N__26708),
            .in1(N__53458),
            .in2(_gnd_net_),
            .in3(N__30682),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNO_0_3_LC_9_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNO_0_3_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNO_0_3_LC_9_6_4 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \phase_controller_inst2.state_RNO_0_3_LC_9_6_4  (
            .in0(N__26752),
            .in1(N__28691),
            .in2(N__26599),
            .in3(N__26575),
            .lcout(\phase_controller_inst2.state_ns_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_LC_9_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_9_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_9_7_2 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_9_7_2  (
            .in0(N__26705),
            .in1(N__26758),
            .in2(N__28699),
            .in3(N__26730),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53839),
            .ce(),
            .sr(N__53340));
    defparam \phase_controller_inst2.state_1_LC_9_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_9_7_3 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \phase_controller_inst2.state_1_LC_9_7_3  (
            .in0(N__26833),
            .in1(N__26786),
            .in2(N__26731),
            .in3(N__26654),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53839),
            .ce(),
            .sr(N__53340));
    defparam \phase_controller_inst2.stoper_hc.running_LC_9_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_9_7_4 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_9_7_4  (
            .in0(N__26704),
            .in1(N__26676),
            .in2(N__30685),
            .in3(N__31122),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53839),
            .ce(),
            .sr(N__53340));
    defparam \phase_controller_inst2.state_2_LC_9_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_9_7_5 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst2.state_2_LC_9_7_5  (
            .in0(N__26759),
            .in1(N__28695),
            .in2(N__26732),
            .in3(N__26653),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53839),
            .ce(),
            .sr(N__53340));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_6  (
            .in0(N__26706),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53839),
            .ce(),
            .sr(N__53340));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_7 .LUT_INIT=16'b1100111000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_7  (
            .in0(N__26677),
            .in1(N__26652),
            .in2(N__31124),
            .in3(N__26660),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53839),
            .ce(),
            .sr(N__53340));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_9_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_9_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33311),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53832),
            .ce(N__37649),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_9_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_9_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_11_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33460),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53832),
            .ce(N__37649),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_9_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_9_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_28_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27794),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53827),
            .ce(N__40966),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_9_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_9_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34307),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53821),
            .ce(N__34247),
            .sr(N__53350));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_9_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_9_11_0 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_9_11_0  (
            .in0(N__29592),
            .in1(N__49118),
            .in2(N__26867),
            .in3(N__26851),
            .lcout(),
            .ltout(\phase_controller_inst1.state_ns_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_9_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_9_11_1 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \phase_controller_inst1.state_3_LC_9_11_1  (
            .in0(N__26980),
            .in1(N__26918),
            .in2(N__26894),
            .in3(N__26891),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53811),
            .ce(),
            .sr(N__53358));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_9_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_9_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_9_11_2  (
            .in0(N__37249),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37276),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un4_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_9_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_9_11_3 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_9_11_3  (
            .in0(N__29019),
            .in1(N__26866),
            .in2(N__26870),
            .in3(N__28369),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53811),
            .ce(),
            .sr(N__53358));
    defparam \phase_controller_inst1.state_0_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_9_11_4 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst1.state_0_LC_9_11_4  (
            .in0(N__26865),
            .in1(N__29614),
            .in2(N__30731),
            .in3(N__26852),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53811),
            .ce(),
            .sr(N__53358));
    defparam \phase_controller_inst1.start_timer_tr_LC_9_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_9_11_5 .LUT_INIT=16'b1011101011111010;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_9_11_5  (
            .in0(N__29756),
            .in1(N__29613),
            .in2(N__37287),
            .in3(N__30729),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53811),
            .ce(),
            .sr(N__53358));
    defparam \phase_controller_inst1.stoper_tr.running_LC_9_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_9_11_7 .LUT_INIT=16'b1111001001110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_9_11_7  (
            .in0(N__37277),
            .in1(N__37250),
            .in2(N__29026),
            .in3(N__28370),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53811),
            .ce(),
            .sr(N__53358));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_9_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_9_12_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_9_12_1  (
            .in0(N__29785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_9_12_4  (
            .in0(N__32552),
            .in1(N__26843),
            .in2(_gnd_net_),
            .in3(N__31734),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(elapsed_time_ns_1_RNIJI91B_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_9_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_9_12_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26837),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_13_0  (
            .in0(N__32638),
            .in1(N__27064),
            .in2(N__32621),
            .in3(N__27073),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_9_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_9_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_9_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34340),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53796),
            .ce(N__34246),
            .sr(N__53368));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_9_13_2  (
            .in0(N__31732),
            .in1(N__27044),
            .in2(_gnd_net_),
            .in3(N__27074),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_13_4  (
            .in0(N__31733),
            .in1(N__27023),
            .in2(_gnd_net_),
            .in3(N__27065),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_9_13_5  (
            .in0(N__31727),
            .in1(N__27053),
            .in2(_gnd_net_),
            .in3(N__32639),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(elapsed_time_ns_1_RNIFE91B_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_9_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_9_13_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27047),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_14_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_14_0  (
            .in0(N__27043),
            .in1(N__41072),
            .in2(N__27032),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__27011),
            .in2(_gnd_net_),
            .in3(N__27022),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__27005),
            .in2(_gnd_net_),
            .in3(N__26999),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__29966),
            .in2(_gnd_net_),
            .in3(N__27224),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__29891),
            .in2(_gnd_net_),
            .in3(N__27203),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__29807),
            .in2(_gnd_net_),
            .in3(N__27182),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__27179),
            .in2(_gnd_net_),
            .in3(N__27149),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__29723),
            .in2(_gnd_net_),
            .in3(N__27128),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__29792),
            .in2(_gnd_net_),
            .in3(N__27113),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__30029),
            .in2(_gnd_net_),
            .in3(N__27098),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__29948),
            .in2(_gnd_net_),
            .in3(N__27077),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__30044),
            .in2(_gnd_net_),
            .in3(N__27413),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__29741),
            .in2(_gnd_net_),
            .in3(N__27389),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__27386),
            .in2(_gnd_net_),
            .in3(N__27356),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_15_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27353),
            .in3(N__27323),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__30062),
            .in2(_gnd_net_),
            .in3(N__27302),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_16_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30014),
            .in3(N__27287),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__30119),
            .in2(_gnd_net_),
            .in3(N__27272),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__30401),
            .in2(_gnd_net_),
            .in3(N__27248),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_16_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29933),
            .in3(N__27611),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__27608),
            .in2(_gnd_net_),
            .in3(N__27578),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__31628),
            .in2(_gnd_net_),
            .in3(N__27557),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__27554),
            .in2(_gnd_net_),
            .in3(N__27530),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__29906),
            .in2(_gnd_net_),
            .in3(N__27509),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__30077),
            .in2(_gnd_net_),
            .in3(N__27494),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__30134),
            .in2(_gnd_net_),
            .in3(N__27479),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__30092),
            .in2(_gnd_net_),
            .in3(N__27458),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__30245),
            .in2(_gnd_net_),
            .in3(N__27854),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__27767),
            .in2(_gnd_net_),
            .in3(N__27830),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__29990),
            .in2(_gnd_net_),
            .in3(N__27809),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_17_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_17_6  (
            .in0(N__27806),
            .in1(N__41074),
            .in2(_gnd_net_),
            .in3(N__27797),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_9_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_9_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30112),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_9_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_9_18_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_9_18_0  (
            .in0(N__27761),
            .in1(N__40985),
            .in2(N__27743),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_0 ),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_9_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_9_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__27734),
            .in2(N__27707),
            .in3(N__27722),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_9_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_9_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__27695),
            .in2(N__27668),
            .in3(N__27683),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_9_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_9_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__27659),
            .in2(N__28112),
            .in3(N__27647),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_9_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_9_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__28103),
            .in2(N__28079),
            .in3(N__28094),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_9_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_9_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_9_18_5  (
            .in0(N__28067),
            .in1(N__28052),
            .in2(N__28043),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_9_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_9_18_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_9_18_6  (
            .in0(N__28034),
            .in1(N__28019),
            .in2(N__28010),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_9_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_9_18_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_9_18_7  (
            .in0(N__28001),
            .in1(N__27983),
            .in2(N__27974),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_9_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_9_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__27932),
            .in2(N__27965),
            .in3(N__27950),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_8 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_9_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_9_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__27926),
            .in2(N__27899),
            .in3(N__27914),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_9_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_9_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__27860),
            .in2(N__27890),
            .in3(N__27875),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_9_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_9_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__28328),
            .in2(N__28301),
            .in3(N__28316),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_9_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_9_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__28262),
            .in2(N__28292),
            .in3(N__28277),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_9_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_9_19_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_9_19_5  (
            .in0(N__28256),
            .in1(N__28241),
            .in2(N__28229),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_9_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_9_19_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_9_19_6  (
            .in0(N__28220),
            .in1(N__28205),
            .in2(N__28193),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_9_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_9_19_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_9_19_7  (
            .in0(N__28184),
            .in1(N__28169),
            .in2(N__28157),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_9_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_9_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__28574),
            .in2(N__28148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_9_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_9_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__28133),
            .in2(N__28124),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_9_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_9_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__30416),
            .in2(N__30170),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_9_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_9_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__28523),
            .in2(N__30302),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_9_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_9_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__28382),
            .in2(N__28853),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_9_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_9_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__28478),
            .in2(N__28394),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_9_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_9_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__28529),
            .in2(N__28337),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_9_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_9_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__29039),
            .in2(N__28928),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_9_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_9_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28373),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_9_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_9_21_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__37242),
            .in2(_gnd_net_),
            .in3(N__28363),
            .lcout(\phase_controller_inst1.stoper_tr.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_9_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_9_21_3 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_9_21_3  (
            .in0(N__28567),
            .in1(N__28967),
            .in2(_gnd_net_),
            .in3(N__28546),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_9_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_9_21_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_9_21_4  (
            .in0(N__28658),
            .in1(N__28638),
            .in2(N__28618),
            .in3(N__28592),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_9_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_9_21_5 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_9_21_5  (
            .in0(N__28568),
            .in1(N__28968),
            .in2(_gnd_net_),
            .in3(N__28547),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_9_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_9_21_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_9_21_6  (
            .in0(N__30385),
            .in1(N__30363),
            .in2(N__30343),
            .in3(N__30316),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_22_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28517),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53757),
            .ce(N__40915),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_22_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28498),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53757),
            .ce(N__40915),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_22_4 .LUT_INIT=16'b0100010011010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_22_4  (
            .in0(N__28450),
            .in1(N__28436),
            .in2(N__28424),
            .in3(N__28408),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28469),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53757),
            .ce(N__40915),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_22_6 .LUT_INIT=16'b1101010011011101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_22_6  (
            .in0(N__28449),
            .in1(N__28435),
            .in2(N__28423),
            .in3(N__28407),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_23_0 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_23_0  (
            .in0(N__28861),
            .in1(N__28878),
            .in2(N__28916),
            .in3(N__28891),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_9_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_9_23_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_9_23_2  (
            .in0(N__28941),
            .in1(N__28986),
            .in2(_gnd_net_),
            .in3(N__28972),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_9_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_9_23_4 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_9_23_4  (
            .in0(N__29030),
            .in1(N__37293),
            .in2(_gnd_net_),
            .in3(N__37238),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_9_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_9_23_5 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_9_23_5  (
            .in0(N__28987),
            .in1(_gnd_net_),
            .in2(N__28973),
            .in3(N__28942),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_23_7 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_23_7  (
            .in0(N__28908),
            .in1(N__28892),
            .in2(N__28880),
            .in3(N__28862),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_9_24_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_9_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37243),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_9_28_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_28_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28706),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53729),
            .ce(),
            .sr(N__53424));
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_10_2_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_10_2_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_10_2_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_0_LC_10_2_0  (
            .in0(N__29348),
            .in1(N__30619),
            .in2(N__30638),
            .in3(N__30637),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_2_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_0 ),
            .clk(N__53851),
            .ce(N__29260),
            .sr(N__53319));
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_10_2_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_10_2_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_10_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_1_LC_10_2_1  (
            .in0(N__29390),
            .in1(N__30598),
            .in2(_gnd_net_),
            .in3(N__28661),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_1 ),
            .clk(N__53851),
            .ce(N__29260),
            .sr(N__53319));
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_10_2_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_10_2_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_10_2_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_2_LC_10_2_2  (
            .in0(N__29349),
            .in1(N__30571),
            .in2(_gnd_net_),
            .in3(N__29066),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_2 ),
            .clk(N__53851),
            .ce(N__29260),
            .sr(N__53319));
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_10_2_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_10_2_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_10_2_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_3_LC_10_2_3  (
            .in0(N__29391),
            .in1(N__30547),
            .in2(_gnd_net_),
            .in3(N__29063),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_3 ),
            .clk(N__53851),
            .ce(N__29260),
            .sr(N__53319));
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_10_2_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_10_2_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_10_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_4_LC_10_2_4  (
            .in0(N__29350),
            .in1(N__30526),
            .in2(_gnd_net_),
            .in3(N__29060),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_4 ),
            .clk(N__53851),
            .ce(N__29260),
            .sr(N__53319));
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_10_2_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_10_2_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_10_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_5_LC_10_2_5  (
            .in0(N__29392),
            .in1(N__30925),
            .in2(_gnd_net_),
            .in3(N__29057),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_5 ),
            .clk(N__53851),
            .ce(N__29260),
            .sr(N__53319));
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_10_2_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_10_2_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_10_2_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_6_LC_10_2_6  (
            .in0(N__29351),
            .in1(N__30904),
            .in2(_gnd_net_),
            .in3(N__29054),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_6 ),
            .clk(N__53851),
            .ce(N__29260),
            .sr(N__53319));
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_10_2_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_10_2_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_10_2_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_7_LC_10_2_7  (
            .in0(N__29393),
            .in1(N__30883),
            .in2(_gnd_net_),
            .in3(N__29051),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_7 ),
            .clk(N__53851),
            .ce(N__29260),
            .sr(N__53319));
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_10_3_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_10_3_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_10_3_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_8_LC_10_3_0  (
            .in0(N__29347),
            .in1(N__30859),
            .in2(_gnd_net_),
            .in3(N__29048),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_10_3_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_8 ),
            .clk(N__53849),
            .ce(N__29256),
            .sr(N__53321));
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_10_3_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_10_3_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_10_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_9_LC_10_3_1  (
            .in0(N__29359),
            .in1(N__30835),
            .in2(_gnd_net_),
            .in3(N__29045),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_9 ),
            .clk(N__53849),
            .ce(N__29256),
            .sr(N__53321));
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_10_3_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_10_3_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_10_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_10_LC_10_3_2  (
            .in0(N__29344),
            .in1(N__30811),
            .in2(_gnd_net_),
            .in3(N__29042),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_10 ),
            .clk(N__53849),
            .ce(N__29256),
            .sr(N__53321));
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_10_3_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_10_3_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_10_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_11_LC_10_3_3  (
            .in0(N__29356),
            .in1(N__30787),
            .in2(_gnd_net_),
            .in3(N__29093),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_11 ),
            .clk(N__53849),
            .ce(N__29256),
            .sr(N__53321));
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_10_3_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_10_3_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_10_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_12_LC_10_3_4  (
            .in0(N__29345),
            .in1(N__30760),
            .in2(_gnd_net_),
            .in3(N__29090),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_12 ),
            .clk(N__53849),
            .ce(N__29256),
            .sr(N__53321));
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_10_3_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_10_3_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_10_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_13_LC_10_3_5  (
            .in0(N__29357),
            .in1(N__31096),
            .in2(_gnd_net_),
            .in3(N__29087),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_13 ),
            .clk(N__53849),
            .ce(N__29256),
            .sr(N__53321));
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_10_3_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_10_3_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_10_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_14_LC_10_3_6  (
            .in0(N__29346),
            .in1(N__31069),
            .in2(_gnd_net_),
            .in3(N__29084),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_14 ),
            .clk(N__53849),
            .ce(N__29256),
            .sr(N__53321));
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_10_3_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_10_3_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_10_3_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_15_LC_10_3_7  (
            .in0(N__29358),
            .in1(N__31045),
            .in2(_gnd_net_),
            .in3(N__29081),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_15 ),
            .clk(N__53849),
            .ce(N__29256),
            .sr(N__53321));
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_10_4_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_10_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_10_4_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_16_LC_10_4_0  (
            .in0(N__29352),
            .in1(N__29682),
            .in2(_gnd_net_),
            .in3(N__29078),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_10_4_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_16 ),
            .clk(N__53845),
            .ce(N__29261),
            .sr(N__53323));
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_10_4_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_10_4_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_10_4_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_17_LC_10_4_1  (
            .in0(N__29386),
            .in1(N__29715),
            .in2(_gnd_net_),
            .in3(N__29075),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_17 ),
            .clk(N__53845),
            .ce(N__29261),
            .sr(N__53323));
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_10_4_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_10_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_10_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_18_LC_10_4_2  (
            .in0(N__29353),
            .in1(N__29490),
            .in2(_gnd_net_),
            .in3(N__29072),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_18 ),
            .clk(N__53845),
            .ce(N__29261),
            .sr(N__53323));
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_10_4_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_10_4_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_10_4_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_19_LC_10_4_3  (
            .in0(N__29387),
            .in1(N__29463),
            .in2(_gnd_net_),
            .in3(N__29069),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_19 ),
            .clk(N__53845),
            .ce(N__29261),
            .sr(N__53323));
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_10_4_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_10_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_10_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_20_LC_10_4_4  (
            .in0(N__29354),
            .in1(N__29136),
            .in2(_gnd_net_),
            .in3(N__29120),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_20 ),
            .clk(N__53845),
            .ce(N__29261),
            .sr(N__53323));
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_10_4_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_10_4_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_10_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_21_LC_10_4_5  (
            .in0(N__29388),
            .in1(N__29160),
            .in2(_gnd_net_),
            .in3(N__29117),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_21 ),
            .clk(N__53845),
            .ce(N__29261),
            .sr(N__53323));
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_10_4_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_10_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_10_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_22_LC_10_4_6  (
            .in0(N__29355),
            .in1(N__29439),
            .in2(_gnd_net_),
            .in3(N__29114),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_22 ),
            .clk(N__53845),
            .ce(N__29261),
            .sr(N__53323));
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_10_4_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_10_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_10_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_23_LC_10_4_7  (
            .in0(N__29389),
            .in1(N__29415),
            .in2(_gnd_net_),
            .in3(N__29111),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_23 ),
            .clk(N__53845),
            .ce(N__29261),
            .sr(N__53323));
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_10_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_10_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_10_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_24_LC_10_5_0  (
            .in0(N__29378),
            .in1(N__29547),
            .in2(_gnd_net_),
            .in3(N__29108),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_10_5_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_24 ),
            .clk(N__53840),
            .ce(N__29249),
            .sr(N__53326));
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_10_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_10_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_10_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_25_LC_10_5_1  (
            .in0(N__29383),
            .in1(N__29565),
            .in2(_gnd_net_),
            .in3(N__29105),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_25 ),
            .clk(N__53840),
            .ce(N__29249),
            .sr(N__53326));
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_10_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_10_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_10_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_26_LC_10_5_2  (
            .in0(N__29379),
            .in1(N__29511),
            .in2(_gnd_net_),
            .in3(N__29102),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_26 ),
            .clk(N__53840),
            .ce(N__29249),
            .sr(N__53326));
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_10_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_10_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_10_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_27_LC_10_5_3  (
            .in0(N__29384),
            .in1(N__29529),
            .in2(_gnd_net_),
            .in3(N__29099),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_27 ),
            .clk(N__53840),
            .ce(N__29249),
            .sr(N__53326));
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_10_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_10_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_10_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_28_LC_10_5_4  (
            .in0(N__29380),
            .in1(N__29225),
            .in2(_gnd_net_),
            .in3(N__29096),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_28 ),
            .clk(N__53840),
            .ce(N__29249),
            .sr(N__53326));
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_10_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_10_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_10_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_29_LC_10_5_5  (
            .in0(N__29385),
            .in1(N__29210),
            .in2(_gnd_net_),
            .in3(N__29399),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_29 ),
            .clk(N__53840),
            .ce(N__29249),
            .sr(N__53326));
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_10_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_10_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_10_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_30_LC_10_5_6  (
            .in0(N__29381),
            .in1(N__29195),
            .in2(_gnd_net_),
            .in3(N__29396),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_29 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_30 ),
            .clk(N__53840),
            .ce(N__29249),
            .sr(N__53326));
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_10_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_10_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_10_5_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_31_LC_10_5_7  (
            .in0(N__29180),
            .in1(N__29382),
            .in2(_gnd_net_),
            .in3(N__29264),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53840),
            .ce(N__29249),
            .sr(N__53326));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_10_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_10_6_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_10_6_0  (
            .in0(N__29224),
            .in1(N__29209),
            .in2(_gnd_net_),
            .in3(N__29649),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_10_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_10_6_1 .LUT_INIT=16'b1011101100101011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_10_6_1  (
            .in0(N__33226),
            .in1(N__29161),
            .in2(N__29143),
            .in3(N__31219),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_10_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_10_6_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_10_6_2  (
            .in0(N__29223),
            .in1(N__29208),
            .in2(_gnd_net_),
            .in3(N__29648),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_10_6_3 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_10_6_3  (
            .in0(N__29650),
            .in1(N__29179),
            .in2(_gnd_net_),
            .in3(N__29193),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_10_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_10_6_4 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_10_6_4  (
            .in0(N__29194),
            .in1(N__29178),
            .in2(_gnd_net_),
            .in3(N__29651),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_10_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_10_6_5 .LUT_INIT=16'b0010101100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_10_6_5  (
            .in0(N__33227),
            .in1(N__29162),
            .in2(N__29144),
            .in3(N__31220),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_10_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_10_6_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_10_6_6  (
            .in0(N__29666),
            .in1(N__29467),
            .in2(N__29495),
            .in3(N__31238),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_10_7_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_10_7_0  (
            .in0(N__31307),
            .in1(N__29567),
            .in2(N__31208),
            .in3(N__29549),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_10_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_10_7_2 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_10_7_2  (
            .in0(N__31306),
            .in1(N__29566),
            .in2(N__31207),
            .in3(N__29548),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_10_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_10_7_4 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_10_7_4  (
            .in0(N__29630),
            .in1(N__29531),
            .in2(N__31190),
            .in3(N__29513),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_10_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_10_7_6 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_10_7_6  (
            .in0(N__29629),
            .in1(N__29530),
            .in2(N__31189),
            .in3(N__29512),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_10_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_10_8_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_10_8_0  (
            .in0(N__29665),
            .in1(N__29491),
            .in2(N__29471),
            .in3(N__31234),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_10_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_10_8_4 .LUT_INIT=16'b0100111100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_10_8_4  (
            .in0(N__29441),
            .in1(N__31247),
            .in2(N__29423),
            .in3(N__31256),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_10_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_10_8_6 .LUT_INIT=16'b1101111100001101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_10_8_6  (
            .in0(N__29440),
            .in1(N__31246),
            .in2(N__29422),
            .in3(N__31255),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_10_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_10_9_0 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_10_9_0  (
            .in0(N__29717),
            .in1(N__29699),
            .in2(N__29690),
            .in3(N__31316),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_10_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_10_9_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_16_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__33982),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53812),
            .ce(N__33374),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_10_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_10_9_2 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_10_9_2  (
            .in0(N__29716),
            .in1(N__29698),
            .in2(N__29689),
            .in3(N__31315),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_10_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_10_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_18_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34642),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53812),
            .ce(N__33374),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_10_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_28_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36482),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53803),
            .ce(N__33375),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_10_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_26_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33686),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53803),
            .ce(N__33375),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_10_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_10_11_0 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.state_1_LC_10_11_0  (
            .in0(N__29773),
            .in1(N__29618),
            .in2(N__34154),
            .in3(N__30722),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53797),
            .ce(),
            .sr(N__53346));
    defparam \phase_controller_inst1.state_2_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_10_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_10_11_1 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_10_11_1  (
            .in0(N__29594),
            .in1(N__29774),
            .in2(N__49129),
            .in3(N__34153),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53797),
            .ce(),
            .sr(N__53346));
    defparam \phase_controller_inst1.start_timer_hc_LC_10_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_10_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_10_11_3 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_10_11_3  (
            .in0(N__29593),
            .in1(N__34022),
            .in2(N__49128),
            .in3(N__29772),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53797),
            .ce(),
            .sr(N__53346));
    defparam \phase_controller_inst1.stoper_hc.running_LC_10_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_10_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_10_11_6 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_10_11_6  (
            .in0(N__34021),
            .in1(N__34198),
            .in2(N__34547),
            .in3(N__34178),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53797),
            .ce(),
            .sr(N__53346));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_10_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_10_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_10_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34023),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53797),
            .ce(),
            .sr(N__53346));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_10_12_0  (
            .in0(N__31759),
            .in1(N__30004),
            .in2(_gnd_net_),
            .in3(N__33143),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_10_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_10_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_10_12_2  (
            .in0(N__31757),
            .in1(N__33011),
            .in2(_gnd_net_),
            .in3(N__29786),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_12_3  (
            .in0(N__29920),
            .in1(N__32936),
            .in2(_gnd_net_),
            .in3(N__31758),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_12_4  (
            .in0(N__29771),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34144),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_12_5  (
            .in0(N__29750),
            .in1(N__32804),
            .in2(_gnd_net_),
            .in3(N__31756),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_10_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_10_12_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29744),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_12_7 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_10_12_7  (
            .in0(N__34197),
            .in1(N__34017),
            .in2(_gnd_net_),
            .in3(N__34527),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_13_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_13_0  (
            .in0(N__32527),
            .in1(N__29732),
            .in2(_gnd_net_),
            .in3(N__31735),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(elapsed_time_ns_1_RNIKJ91B_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_13_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29726),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_i_LC_10_13_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_i_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_i_LC_10_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un3_threshold_i_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29878),
            .lcout(\pwm_generator_inst.un3_threshold_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_13_3  (
            .in0(N__31736),
            .in1(N__29960),
            .in2(_gnd_net_),
            .in3(N__32849),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_13_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_13_4  (
            .in0(N__32548),
            .in1(N__29828),
            .in2(N__32528),
            .in3(N__30158),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_13_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_13_5  (
            .in0(N__33112),
            .in1(N__30143),
            .in2(N__29822),
            .in3(N__30284),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_13_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__29816),
            .in2(N__29819),
            .in3(N__32573),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(elapsed_time_ns_1_RNIIH91B_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29810),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_14_0  (
            .in0(N__31729),
            .in1(N__29801),
            .in2(_gnd_net_),
            .in3(N__32507),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(elapsed_time_ns_1_RNILK91B_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_10_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_10_14_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29795),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_14_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_10_14_2  (
            .in0(N__31730),
            .in1(N__30056),
            .in2(_gnd_net_),
            .in3(N__32825),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_14_3  (
            .in0(N__32617),
            .in1(N__29975),
            .in2(_gnd_net_),
            .in3(N__31728),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(elapsed_time_ns_1_RNIGF91B_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_14_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29969),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_14_5  (
            .in0(N__29959),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_14_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_14_6  (
            .in0(N__31731),
            .in1(N__29942),
            .in2(_gnd_net_),
            .in3(N__33035),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29936),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_15_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_15_0  (
            .in0(N__29921),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_10_15_1  (
            .in0(N__29900),
            .in1(N__32594),
            .in2(_gnd_net_),
            .in3(N__31766),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(elapsed_time_ns_1_RNIHG91B_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_10_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_10_15_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29894),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_15_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_15_3  (
            .in0(N__29885),
            .in1(N__32729),
            .in2(_gnd_net_),
            .in3(N__31768),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_10_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_10_15_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30065),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_10_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_10_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_10_15_5  (
            .in0(N__30055),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_10_15_6  (
            .in0(N__31767),
            .in1(N__30038),
            .in2(_gnd_net_),
            .in3(N__32870),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_10_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_10_15_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30032),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_16_1  (
            .in0(N__30023),
            .in1(N__32705),
            .in2(_gnd_net_),
            .in3(N__31769),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(elapsed_time_ns_1_RNI4EOBB_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_16_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30017),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_10_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_10_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30005),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_16_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_16_4  (
            .in0(N__31771),
            .in1(N__29984),
            .in2(_gnd_net_),
            .in3(N__32891),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_10_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_10_16_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29978),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_16_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_10_16_6  (
            .in0(N__31770),
            .in1(N__30128),
            .in2(_gnd_net_),
            .in3(N__33068),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_10_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_10_16_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30122),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_17_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_10_17_0  (
            .in0(N__30113),
            .in1(N__33164),
            .in2(_gnd_net_),
            .in3(N__31781),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_10_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_10_17_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_10_17_1  (
            .in0(N__31779),
            .in1(N__30101),
            .in2(_gnd_net_),
            .in3(N__33209),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_10_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_10_17_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30095),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_17_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_17_4  (
            .in0(N__30086),
            .in1(N__31778),
            .in2(_gnd_net_),
            .in3(N__32912),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(elapsed_time_ns_1_RNI3EPBB_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_17_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30080),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_17_6  (
            .in0(N__30071),
            .in1(N__33188),
            .in2(_gnd_net_),
            .in3(N__31780),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_10_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_10_17_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30248),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_10_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_10_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_20_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30239),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53768),
            .ce(N__40941),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_10_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_10_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_21_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30223),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53768),
            .ce(N__40941),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_10_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_10_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_22_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30206),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53768),
            .ce(N__40941),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_10_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_10_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_23_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30184),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53768),
            .ce(N__40941),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_10_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_10_19_0 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_10_19_0  (
            .in0(N__30487),
            .in1(N__30457),
            .in2(N__30443),
            .in3(N__30499),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_10_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_10_19_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__32566),
            .in2(_gnd_net_),
            .in3(N__32587),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_20_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_10_20_3  (
            .in0(N__32839),
            .in1(N__32863),
            .in2(N__32503),
            .in3(N__32818),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_10_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_10_20_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__32767),
            .in2(N__30146),
            .in3(N__32791),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_10_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_10_20_7 .LUT_INIT=16'b0010001010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_10_20_7  (
            .in0(N__30503),
            .in1(N__30488),
            .in2(N__30461),
            .in3(N__30442),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_21_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_10_21_1  (
            .in0(N__30410),
            .in1(N__33047),
            .in2(_gnd_net_),
            .in3(N__31786),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_10_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_10_21_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30404),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_10_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_10_21_3 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_10_21_3  (
            .in0(N__30386),
            .in1(N__30371),
            .in2(N__30347),
            .in3(N__30317),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_10_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_10_21_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_10_21_4  (
            .in0(N__32698),
            .in1(N__32743),
            .in2(N__32725),
            .in3(N__33061),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_10_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_10_21_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_10_21_5  (
            .in0(N__33001),
            .in1(N__33025),
            .in2(N__32983),
            .in3(N__33046),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_10_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_10_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_10_21_6  (
            .in0(N__30293),
            .in1(N__30737),
            .in2(N__30287),
            .in3(N__30254),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_22_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__30272),
            .in2(_gnd_net_),
            .in3(N__35980),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_22_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_10_22_2  (
            .in0(N__33202),
            .in1(N__32884),
            .in2(N__33184),
            .in3(N__32905),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_10_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_10_22_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_10_22_4  (
            .in0(N__33157),
            .in1(N__32950),
            .in2(N__32932),
            .in3(N__33133),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_10_28_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_10_28_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_10_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_10_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30730),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53727),
            .ce(),
            .sr(N__53422));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_3_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_3_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_3_6  (
            .in0(_gnd_net_),
            .in1(N__30686),
            .in2(_gnd_net_),
            .in3(N__31123),
            .lcout(\phase_controller_inst2.stoper_hc.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_4_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__30605),
            .in2(N__33404),
            .in3(N__30623),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_0 ),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_4_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__33083),
            .in2(N__30584),
            .in3(N__30599),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_4_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_4_2  (
            .in0(_gnd_net_),
            .in1(N__33089),
            .in2(N__30557),
            .in3(N__30575),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_4_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(N__30533),
            .in2(N__33242),
            .in3(N__30548),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_4_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_4_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_4_4  (
            .in0(N__30527),
            .in1(N__33266),
            .in2(N__30512),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_4_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_4_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_4_5  (
            .in0(N__30926),
            .in1(N__30911),
            .in2(N__33077),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_4_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_4_6  (
            .in0(_gnd_net_),
            .in1(N__30890),
            .in2(N__33251),
            .in3(N__30905),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_4_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_4_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_4_7  (
            .in0(N__30884),
            .in1(N__30869),
            .in2(N__33260),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_5_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_5_0  (
            .in0(N__30863),
            .in1(N__33410),
            .in2(N__30845),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_8 ),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__30821),
            .in2(N__33275),
            .in3(N__30836),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__33233),
            .in2(N__30797),
            .in3(N__30815),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__33281),
            .in2(N__30773),
            .in3(N__30788),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_5_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_5_4  (
            .in0(N__30761),
            .in1(N__33215),
            .in2(N__30746),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_5_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_5_5  (
            .in0(N__31097),
            .in1(N__33416),
            .in2(N__31082),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(N__33422),
            .in2(N__31055),
            .in3(N__31070),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_5_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_5_7  (
            .in0(N__31046),
            .in1(N__31031),
            .in2(N__33389),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__31025),
            .in2(N__31013),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__30998),
            .in2(N__30992),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__30977),
            .in2(N__30971),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__30962),
            .in2(N__30953),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__30941),
            .in2(N__30935),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__31172),
            .in2(N__31166),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__31157),
            .in2(N__31151),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__31142),
            .in2(N__31136),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31127),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_11_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_11_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_15_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33586),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53813),
            .ce(N__37647),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_11_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_11_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_8_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33496),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53813),
            .ce(N__37647),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_11_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_11_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_5_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33520),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53813),
            .ce(N__37647),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_11_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_11_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_9_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33478),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53813),
            .ce(N__37647),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_11_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_11_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_12_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33436),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53813),
            .ce(N__37647),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_11_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_11_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_14_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33604),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53813),
            .ce(N__37647),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_11_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_11_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_13_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33622),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53813),
            .ce(N__37647),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_11_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_11_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_23_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33719),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53813),
            .ce(N__37647),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_11_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_11_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_23_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33718),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53804),
            .ce(N__33380),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_11_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_22_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33733),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53804),
            .ce(N__33380),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_11_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_11_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_19_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33844),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53804),
            .ce(N__33380),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_11_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_11_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_20_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33559),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53804),
            .ce(N__33380),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_11_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_11_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_25_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33755),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53804),
            .ce(N__33380),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_11_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_27_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33668),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53804),
            .ce(N__33380),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_11_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_11_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_17_LC_11_9_6  (
            .in0(N__34669),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53804),
            .ce(N__33380),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_11_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_11_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_24_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33704),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53804),
            .ce(N__33380),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_10_0 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_10_0  (
            .in0(N__32180),
            .in1(N__31295),
            .in2(N__32210),
            .in3(N__31286),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_11_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_11_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_20_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33560),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53798),
            .ce(N__37635),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_11_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_11_10_2 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_11_10_2  (
            .in0(N__32179),
            .in1(N__31294),
            .in2(N__32209),
            .in3(N__31285),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_11_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_11_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_21_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33541),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53798),
            .ce(N__37635),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_10_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_10_4  (
            .in0(N__31277),
            .in1(N__32453),
            .in2(N__32483),
            .in3(N__31268),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_11_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_11_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_22_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33734),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53798),
            .ce(N__37635),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_11_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_11_10_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_11_10_6  (
            .in0(N__31276),
            .in1(N__32452),
            .in2(N__32482),
            .in3(N__31267),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_11_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_11_11_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_11_11_0  (
            .in0(N__31382),
            .in1(N__32399),
            .in2(N__32428),
            .in3(N__33743),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_11_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_11_11_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_24_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__33703),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53789),
            .ce(N__37642),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_11_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_11_11_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_11_11_2  (
            .in0(N__31381),
            .in1(N__32398),
            .in2(N__32429),
            .in3(N__33742),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_11_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_11_11_4 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_11_11_4  (
            .in0(N__32348),
            .in1(N__31373),
            .in2(N__32375),
            .in3(N__31364),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_11_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_26_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33685),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53789),
            .ce(N__37642),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_11_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_11_11_6 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_11_11_6  (
            .in0(N__32347),
            .in1(N__31372),
            .in2(N__32374),
            .in3(N__31363),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_11_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_27_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33667),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53789),
            .ce(N__37642),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_11_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_11_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__37658),
            .in2(N__31355),
            .in3(N__31964),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_0 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_11_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_11_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__31331),
            .in2(N__31346),
            .in3(N__31946),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_11_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_11_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__33881),
            .in2(N__31325),
            .in3(N__31925),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_11_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_11_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__33815),
            .in2(N__31487),
            .in3(N__31904),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_11_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_11_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__33632),
            .in2(N__31475),
            .in3(N__31883),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_11_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_11_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_11_12_5  (
            .in0(N__32153),
            .in1(N__31463),
            .in2(N__31451),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_11_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_11_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__31439),
            .in2(N__33857),
            .in3(N__32135),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_11_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_11_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_11_12_7  (
            .in0(N__32114),
            .in1(N__31433),
            .in2(N__33791),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_11_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_11_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_11_13_0  (
            .in0(N__32096),
            .in1(N__31427),
            .in2(N__31418),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_8 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_11_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_11_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__31409),
            .in2(N__31400),
            .in3(N__32078),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_11_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_11_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__33764),
            .in2(N__31391),
            .in3(N__32060),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_11_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_11_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__31598),
            .in2(N__31616),
            .in3(N__32039),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_11_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_11_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__31592),
            .in2(N__31580),
            .in3(N__32021),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_11_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_11_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__31571),
            .in2(N__31562),
            .in3(N__32279),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_11_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_11_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_11_13_6  (
            .in0(N__32258),
            .in1(N__31550),
            .in2(N__31538),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_11_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_11_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_11_13_7  (
            .in0(N__32240),
            .in1(N__31514),
            .in2(N__31526),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_11_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_11_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__33989),
            .in2(N__33908),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_11_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_11_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__34649),
            .in2(N__34556),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_11_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_11_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__31508),
            .in2(N__31499),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_11_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_11_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__31862),
            .in2(N__31850),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_11_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_11_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__31835),
            .in2(N__31826),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_11_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_11_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__31814),
            .in2(N__31802),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_11_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_11_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__31985),
            .in2(N__32000),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_11_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_11_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__31991),
            .in2(N__36383),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31790),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_11_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_11_15_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_11_15_2  (
            .in0(N__31637),
            .in1(N__32987),
            .in2(_gnd_net_),
            .in3(N__31785),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_11_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_11_15_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31631),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_11_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_11_15_4 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_11_15_4  (
            .in0(N__32303),
            .in1(N__36405),
            .in2(_gnd_net_),
            .in3(N__32326),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_11_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_11_15_5 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_11_15_5  (
            .in0(N__36407),
            .in1(N__36460),
            .in2(_gnd_net_),
            .in3(N__36430),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_11_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_11_15_6 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_11_15_6  (
            .in0(N__32302),
            .in1(N__36406),
            .in2(_gnd_net_),
            .in3(N__32327),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_11_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_11_15_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__34543),
            .in2(_gnd_net_),
            .in3(N__34167),
            .lcout(\phase_controller_inst1.stoper_hc.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_11_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_11_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_11_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_0_LC_11_16_0  (
            .in0(N__34493),
            .in1(N__31960),
            .in2(N__31979),
            .in3(N__31978),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_0 ),
            .clk(N__53775),
            .ce(N__32676),
            .sr(N__53369));
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_11_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_11_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_11_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_1_LC_11_16_1  (
            .in0(N__34406),
            .in1(N__31942),
            .in2(_gnd_net_),
            .in3(N__31928),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_1 ),
            .clk(N__53775),
            .ce(N__32676),
            .sr(N__53369));
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_11_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_11_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_11_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_2_LC_11_16_2  (
            .in0(N__34494),
            .in1(N__31921),
            .in2(_gnd_net_),
            .in3(N__31907),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_2 ),
            .clk(N__53775),
            .ce(N__32676),
            .sr(N__53369));
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_11_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_11_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_11_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_3_LC_11_16_3  (
            .in0(N__34407),
            .in1(N__31903),
            .in2(_gnd_net_),
            .in3(N__31886),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_3 ),
            .clk(N__53775),
            .ce(N__32676),
            .sr(N__53369));
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_11_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_11_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_11_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_4_LC_11_16_4  (
            .in0(N__34495),
            .in1(N__31879),
            .in2(_gnd_net_),
            .in3(N__31865),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_4 ),
            .clk(N__53775),
            .ce(N__32676),
            .sr(N__53369));
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_11_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_11_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_11_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_5_LC_11_16_5  (
            .in0(N__34408),
            .in1(N__32152),
            .in2(_gnd_net_),
            .in3(N__32138),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_5 ),
            .clk(N__53775),
            .ce(N__32676),
            .sr(N__53369));
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_11_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_11_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_11_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_6_LC_11_16_6  (
            .in0(N__34496),
            .in1(N__32131),
            .in2(_gnd_net_),
            .in3(N__32117),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_6 ),
            .clk(N__53775),
            .ce(N__32676),
            .sr(N__53369));
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_11_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_11_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_11_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_7_LC_11_16_7  (
            .in0(N__34409),
            .in1(N__32113),
            .in2(_gnd_net_),
            .in3(N__32099),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_7 ),
            .clk(N__53775),
            .ce(N__32676),
            .sr(N__53369));
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_11_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_11_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_11_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_8_LC_11_17_0  (
            .in0(N__34436),
            .in1(N__32095),
            .in2(_gnd_net_),
            .in3(N__32081),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_8 ),
            .clk(N__53769),
            .ce(N__32678),
            .sr(N__53373));
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_11_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_11_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_11_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_9_LC_11_17_1  (
            .in0(N__34492),
            .in1(N__32077),
            .in2(_gnd_net_),
            .in3(N__32063),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_9 ),
            .clk(N__53769),
            .ce(N__32678),
            .sr(N__53373));
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_11_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_11_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_10_LC_11_17_2  (
            .in0(N__34433),
            .in1(N__32056),
            .in2(_gnd_net_),
            .in3(N__32042),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_10 ),
            .clk(N__53769),
            .ce(N__32678),
            .sr(N__53373));
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_11_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_11_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_11_LC_11_17_3  (
            .in0(N__34489),
            .in1(N__32038),
            .in2(_gnd_net_),
            .in3(N__32024),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_11 ),
            .clk(N__53769),
            .ce(N__32678),
            .sr(N__53373));
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_11_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_11_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_11_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_12_LC_11_17_4  (
            .in0(N__34434),
            .in1(N__32017),
            .in2(_gnd_net_),
            .in3(N__32003),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_12 ),
            .clk(N__53769),
            .ce(N__32678),
            .sr(N__53373));
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_11_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_11_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_11_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_13_LC_11_17_5  (
            .in0(N__34490),
            .in1(N__32275),
            .in2(_gnd_net_),
            .in3(N__32261),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_13 ),
            .clk(N__53769),
            .ce(N__32678),
            .sr(N__53373));
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_11_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_11_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_11_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_14_LC_11_17_6  (
            .in0(N__34435),
            .in1(N__32257),
            .in2(_gnd_net_),
            .in3(N__32243),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_14 ),
            .clk(N__53769),
            .ce(N__32678),
            .sr(N__53373));
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_11_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_11_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_11_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_15_LC_11_17_7  (
            .in0(N__34491),
            .in1(N__32239),
            .in2(_gnd_net_),
            .in3(N__32225),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_15 ),
            .clk(N__53769),
            .ce(N__32678),
            .sr(N__53373));
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_11_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_11_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_11_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_16_LC_11_18_0  (
            .in0(N__34481),
            .in1(N__33922),
            .in2(_gnd_net_),
            .in3(N__32222),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_16 ),
            .clk(N__53764),
            .ce(N__32677),
            .sr(N__53378));
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_11_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_11_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_11_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_17_LC_11_18_1  (
            .in0(N__34485),
            .in1(N__33949),
            .in2(_gnd_net_),
            .in3(N__32219),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_17 ),
            .clk(N__53764),
            .ce(N__32677),
            .sr(N__53378));
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_11_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_11_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_11_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_18_LC_11_18_2  (
            .in0(N__34482),
            .in1(N__34570),
            .in2(_gnd_net_),
            .in3(N__32216),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_18 ),
            .clk(N__53764),
            .ce(N__32677),
            .sr(N__53378));
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_11_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_11_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_11_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_19_LC_11_18_3  (
            .in0(N__34486),
            .in1(N__34591),
            .in2(_gnd_net_),
            .in3(N__32213),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_19 ),
            .clk(N__53764),
            .ce(N__32677),
            .sr(N__53378));
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_11_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_11_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_11_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_20_LC_11_18_4  (
            .in0(N__34483),
            .in1(N__32197),
            .in2(_gnd_net_),
            .in3(N__32183),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_20 ),
            .clk(N__53764),
            .ce(N__32677),
            .sr(N__53378));
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_11_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_11_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_11_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_21_LC_11_18_5  (
            .in0(N__34487),
            .in1(N__32170),
            .in2(_gnd_net_),
            .in3(N__32156),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_21 ),
            .clk(N__53764),
            .ce(N__32677),
            .sr(N__53378));
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_11_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_11_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_11_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_22_LC_11_18_6  (
            .in0(N__34484),
            .in1(N__32470),
            .in2(_gnd_net_),
            .in3(N__32456),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_22 ),
            .clk(N__53764),
            .ce(N__32677),
            .sr(N__53378));
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_11_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_11_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_11_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_23_LC_11_18_7  (
            .in0(N__34488),
            .in1(N__32446),
            .in2(_gnd_net_),
            .in3(N__32432),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_23 ),
            .clk(N__53764),
            .ce(N__32677),
            .sr(N__53378));
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_11_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_11_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_11_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_24_LC_11_19_0  (
            .in0(N__34455),
            .in1(N__32416),
            .in2(_gnd_net_),
            .in3(N__32402),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_24 ),
            .clk(N__53758),
            .ce(N__32675),
            .sr(N__53384));
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_11_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_11_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_11_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_25_LC_11_19_1  (
            .in0(N__34460),
            .in1(N__32392),
            .in2(_gnd_net_),
            .in3(N__32378),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_25 ),
            .clk(N__53758),
            .ce(N__32675),
            .sr(N__53384));
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_11_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_11_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_11_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_26_LC_11_19_2  (
            .in0(N__34456),
            .in1(N__32367),
            .in2(_gnd_net_),
            .in3(N__32351),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_26 ),
            .clk(N__53758),
            .ce(N__32675),
            .sr(N__53384));
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_11_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_11_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_11_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_27_LC_11_19_3  (
            .in0(N__34461),
            .in1(N__32346),
            .in2(_gnd_net_),
            .in3(N__32330),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_27 ),
            .clk(N__53758),
            .ce(N__32675),
            .sr(N__53384));
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_11_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_11_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_11_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_28_LC_11_19_4  (
            .in0(N__34457),
            .in1(N__32320),
            .in2(_gnd_net_),
            .in3(N__32306),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_28 ),
            .clk(N__53758),
            .ce(N__32675),
            .sr(N__53384));
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_11_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_11_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_11_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_29_LC_11_19_5  (
            .in0(N__34462),
            .in1(N__32296),
            .in2(_gnd_net_),
            .in3(N__32282),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_29 ),
            .clk(N__53758),
            .ce(N__32675),
            .sr(N__53384));
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_11_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_11_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_11_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_30_LC_11_19_6  (
            .in0(N__34458),
            .in1(N__36429),
            .in2(_gnd_net_),
            .in3(N__32684),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_30 ),
            .clk(N__53758),
            .ce(N__32675),
            .sr(N__53384));
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_11_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_11_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_11_19_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_31_LC_11_19_7  (
            .in0(N__36456),
            .in1(N__34459),
            .in2(_gnd_net_),
            .in3(N__32681),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53758),
            .ce(N__32675),
            .sr(N__53384));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_11_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_11_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_11_20_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__34881),
            .in2(N__34333),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__53752),
            .ce(N__34259),
            .sr(N__53390));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_11_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_11_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_11_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__34860),
            .in2(N__34297),
            .in3(N__32597),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__53752),
            .ce(N__34259),
            .sr(N__53390));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_11_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_11_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_11_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__34882),
            .in2(N__34840),
            .in3(N__32576),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__53752),
            .ce(N__34259),
            .sr(N__53390));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_11_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_11_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_11_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__34812),
            .in2(N__34865),
            .in3(N__32555),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__53752),
            .ce(N__34259),
            .sr(N__53390));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_11_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_11_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_11_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(N__34788),
            .in2(N__34841),
            .in3(N__32531),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__53752),
            .ce(N__34259),
            .sr(N__53390));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_11_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_11_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_11_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__34764),
            .in2(N__34817),
            .in3(N__32510),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__53752),
            .ce(N__34259),
            .sr(N__53390));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_11_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_11_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_11_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__34740),
            .in2(N__34793),
            .in3(N__32486),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__53752),
            .ce(N__34259),
            .sr(N__53390));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_11_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_11_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_11_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(N__34716),
            .in2(N__34769),
            .in3(N__32852),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__53752),
            .ce(N__34259),
            .sr(N__53390));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_11_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_11_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_11_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__34692),
            .in2(N__34745),
            .in3(N__32828),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__53747),
            .ce(N__34269),
            .sr(N__53400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_11_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_11_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_11_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__35070),
            .in2(N__34721),
            .in3(N__32807),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__53747),
            .ce(N__34269),
            .sr(N__53400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_11_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_11_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_11_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__35046),
            .in2(N__34697),
            .in3(N__32780),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__53747),
            .ce(N__34269),
            .sr(N__53400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_11_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_11_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_11_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__35022),
            .in2(N__35075),
            .in3(N__32756),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__53747),
            .ce(N__34269),
            .sr(N__53400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_11_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_11_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_11_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__34998),
            .in2(N__35051),
            .in3(N__32732),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__53747),
            .ce(N__34269),
            .sr(N__53400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_11_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_11_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_11_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(N__34974),
            .in2(N__35027),
            .in3(N__32708),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__53747),
            .ce(N__34269),
            .sr(N__53400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_11_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_11_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_11_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__34950),
            .in2(N__35003),
            .in3(N__32687),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__53747),
            .ce(N__34269),
            .sr(N__53400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_11_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_11_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_11_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__34926),
            .in2(N__34979),
            .in3(N__33050),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__53747),
            .ce(N__34269),
            .sr(N__53400));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_11_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_11_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_11_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__34902),
            .in2(N__34955),
            .in3(N__33038),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__53742),
            .ce(N__34271),
            .sr(N__53406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_11_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_11_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_11_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__35256),
            .in2(N__34931),
            .in3(N__33014),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__53742),
            .ce(N__34271),
            .sr(N__53406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_11_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_11_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_11_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__35232),
            .in2(N__34907),
            .in3(N__32990),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__53742),
            .ce(N__34271),
            .sr(N__53406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_11_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_11_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_11_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__35208),
            .in2(N__35261),
            .in3(N__32966),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__53742),
            .ce(N__34271),
            .sr(N__53406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_11_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_11_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_11_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__35184),
            .in2(N__35237),
            .in3(N__32939),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__53742),
            .ce(N__34271),
            .sr(N__53406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_11_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_11_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_11_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__35160),
            .in2(N__35213),
            .in3(N__32915),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__53742),
            .ce(N__34271),
            .sr(N__53406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_11_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_11_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_11_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__35136),
            .in2(N__35189),
            .in3(N__32894),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__53742),
            .ce(N__34271),
            .sr(N__53406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_11_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_11_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_11_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__35112),
            .in2(N__35165),
            .in3(N__32873),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__53742),
            .ce(N__34271),
            .sr(N__53406));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_11_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_11_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_11_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__35091),
            .in2(N__35141),
            .in3(N__33191),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__53737),
            .ce(N__34270),
            .sr(N__53410));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_11_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_11_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_11_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__35661),
            .in2(N__35117),
            .in3(N__33167),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__53737),
            .ce(N__34270),
            .sr(N__53410));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_11_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_11_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_11_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__35092),
            .in2(N__35642),
            .in3(N__33146),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__53737),
            .ce(N__34270),
            .sr(N__53410));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_11_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_11_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_11_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(N__35494),
            .in2(N__35666),
            .in3(N__33122),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__53737),
            .ce(N__34270),
            .sr(N__53410));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_11_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_11_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_11_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33119),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53737),
            .ce(N__34270),
            .sr(N__53410));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33895),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53833),
            .ce(N__33367),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33307),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53833),
            .ce(N__33367),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33524),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53833),
            .ce(N__33367),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33461),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53828),
            .ce(N__33352),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33482),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53828),
            .ce(N__33352),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33649),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53828),
            .ce(N__33352),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33808),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53828),
            .ce(N__33352),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33874),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53828),
            .ce(N__33352),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33829),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53828),
            .ce(N__33352),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33781),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53822),
            .ce(N__33376),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33545),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53822),
            .ce(N__33376),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33440),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53822),
            .ce(N__33376),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33608),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53822),
            .ce(N__33376),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33626),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53822),
            .ce(N__33376),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33500),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53822),
            .ce(N__33376),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_12_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_12_6_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_0_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__37735),
            .in2(_gnd_net_),
            .in3(N__37680),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53822),
            .ce(N__33376),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33590),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53822),
            .ce(N__33376),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_12_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_12_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__33317),
            .in2(N__37681),
            .in3(N__37719),
            .lcout(\phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ),
            .ltout(),
            .carryin(bfn_12_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_12_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_12_7_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_12_7_1  (
            .in0(N__36086),
            .in1(N__36085),
            .in2(N__42772),
            .in3(N__33290),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_1),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_12_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_12_7_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_12_7_2  (
            .in0(N__36065),
            .in1(N__36064),
            .in2(N__42776),
            .in3(N__33287),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_2),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_12_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_12_7_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_12_7_3  (
            .in0(N__36050),
            .in1(N__36049),
            .in2(N__42773),
            .in3(N__33284),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_3),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_12_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_12_7_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_12_7_4  (
            .in0(N__36035),
            .in1(N__36034),
            .in2(N__42777),
            .in3(N__33527),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_4),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_12_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_12_7_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_12_7_5  (
            .in0(N__36020),
            .in1(N__36019),
            .in2(N__42774),
            .in3(N__33509),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_5),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_12_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_12_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_12_7_6  (
            .in0(N__36005),
            .in1(N__36004),
            .in2(N__42778),
            .in3(N__33506),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_6),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_12_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_12_7_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_12_7_7  (
            .in0(N__36239),
            .in1(N__36238),
            .in2(N__42775),
            .in3(N__33503),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_7),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_12_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_12_8_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_12_8_0  (
            .in0(N__36224),
            .in1(N__36223),
            .in2(N__42770),
            .in3(N__33485),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_8),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_12_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_12_8_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_12_8_1  (
            .in0(N__36209),
            .in1(N__36208),
            .in2(N__42767),
            .in3(N__33467),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_9),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_12_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_12_8_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_12_8_2  (
            .in0(N__36194),
            .in1(N__36193),
            .in2(N__42771),
            .in3(N__33464),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_10),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_12_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_12_8_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_12_8_3  (
            .in0(N__36179),
            .in1(N__36178),
            .in2(N__42764),
            .in3(N__33443),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_11),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_12_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_12_8_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_12_8_4  (
            .in0(N__36155),
            .in1(N__36154),
            .in2(N__42768),
            .in3(N__33425),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_12),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_12_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_12_8_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_12_8_5  (
            .in0(N__36140),
            .in1(N__36139),
            .in2(N__42765),
            .in3(N__33611),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_13),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_12_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_12_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_12_8_6  (
            .in0(N__36125),
            .in1(N__36124),
            .in2(N__42769),
            .in3(N__33593),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_14),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_12_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_12_8_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_12_8_7  (
            .in0(N__36110),
            .in1(N__36109),
            .in2(N__42766),
            .in3(N__33575),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_15),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_12_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_12_9_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_12_9_0  (
            .in0(N__36368),
            .in1(N__36367),
            .in2(N__42705),
            .in3(N__33572),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_16),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_12_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_12_9_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_12_9_1  (
            .in0(N__36353),
            .in1(N__36352),
            .in2(N__42709),
            .in3(N__33569),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_17),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_12_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_12_9_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_12_9_2  (
            .in0(N__36338),
            .in1(N__36337),
            .in2(N__42706),
            .in3(N__33566),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_18),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_12_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_12_9_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_12_9_3  (
            .in0(N__36314),
            .in1(N__36313),
            .in2(N__42710),
            .in3(N__33563),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_19),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_12_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_12_9_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_12_9_4  (
            .in0(N__36299),
            .in1(N__36298),
            .in2(N__42707),
            .in3(N__33548),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_20),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_12_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_12_9_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_12_9_5  (
            .in0(N__36284),
            .in1(N__36283),
            .in2(N__42711),
            .in3(N__33530),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_21),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_12_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_12_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_12_9_6  (
            .in0(N__36269),
            .in1(N__36268),
            .in2(N__42708),
            .in3(N__33722),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_22),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_12_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_12_9_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_12_9_7  (
            .in0(N__36254),
            .in1(N__36253),
            .in2(N__42712),
            .in3(N__33707),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_23),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_12_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_12_10_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_12_10_0  (
            .in0(N__36557),
            .in1(N__36556),
            .in2(N__42630),
            .in3(N__33692),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_24),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_12_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_12_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_12_10_1  (
            .in0(N__36542),
            .in1(N__36541),
            .in2(N__42632),
            .in3(N__33689),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_25),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_12_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_12_10_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_12_10_2  (
            .in0(N__36527),
            .in1(N__36526),
            .in2(N__42631),
            .in3(N__33671),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_26),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_12_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_12_10_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_12_10_3  (
            .in0(N__36512),
            .in1(N__36511),
            .in2(N__42633),
            .in3(N__33656),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_27),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_12_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_12_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33653),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_12_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_12_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_4_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33650),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53787),
            .ce(N__37622),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_12_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_2_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33899),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53787),
            .ce(N__37622),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_12_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_6_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33875),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53787),
            .ce(N__37622),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_12_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_12_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_19_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33848),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53787),
            .ce(N__37622),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_12_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_12_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_3_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33833),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53787),
            .ce(N__37622),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_12_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_12_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_7_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33809),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53787),
            .ce(N__37622),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_12_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_12_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_10_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33782),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53787),
            .ce(N__37622),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_12_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_12_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_25_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33754),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53787),
            .ce(N__37622),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_0 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_0  (
            .in0(N__34359),
            .in1(_gnd_net_),
            .in2(N__48854),
            .in3(N__48877),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_168_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_12_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_12_12_1  (
            .in0(N__48878),
            .in1(N__34360),
            .in2(_gnd_net_),
            .in3(N__48853),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53784),
            .ce(),
            .sr(N__53341));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__34358),
            .in2(_gnd_net_),
            .in3(N__48849),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_167_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_12_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_12_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__34030),
            .in2(_gnd_net_),
            .in3(N__34546),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un4_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_12_6 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_12_12_6  (
            .in0(N__34205),
            .in1(N__34143),
            .in2(N__34181),
            .in3(N__34174),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53784),
            .ce(),
            .sr(N__53341));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_12_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_12_13_0 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_12_13_0  (
            .in0(N__34123),
            .in1(N__34093),
            .in2(_gnd_net_),
            .in3(N__34070),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_12_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_12_13_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_12_13_3  (
            .in0(N__34031),
            .in1(N__53459),
            .in2(_gnd_net_),
            .in3(N__34545),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_13_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_12_13_7  (
            .in0(N__49943),
            .in1(N__39049),
            .in2(N__49756),
            .in3(N__39011),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_14_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_14_0  (
            .in0(N__33965),
            .in1(N__33956),
            .in2(N__33935),
            .in3(N__34658),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_12_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_16_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33983),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53779),
            .ce(N__37600),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_12_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_12_14_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_12_14_2  (
            .in0(N__33964),
            .in1(N__33955),
            .in2(N__33934),
            .in3(N__34657),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_12_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_12_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_17_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34673),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53779),
            .ce(N__37600),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_12_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_12_14_4 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_12_14_4  (
            .in0(N__34625),
            .in1(N__34616),
            .in2(N__34603),
            .in3(N__34577),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_12_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_12_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_18_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34643),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53779),
            .ce(N__37600),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_12_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_12_14_6 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_12_14_6  (
            .in0(N__34624),
            .in1(N__34615),
            .in2(N__34604),
            .in3(N__34576),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_12_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_12_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34544),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34361),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_12_19_0  (
            .in0(N__35586),
            .in1(N__34326),
            .in2(_gnd_net_),
            .in3(N__34310),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__53751),
            .ce(N__35458),
            .sr(N__53379));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_12_19_1  (
            .in0(N__35621),
            .in1(N__34290),
            .in2(_gnd_net_),
            .in3(N__34274),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__53751),
            .ce(N__35458),
            .sr(N__53379));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_12_19_2  (
            .in0(N__35587),
            .in1(N__34883),
            .in2(_gnd_net_),
            .in3(N__34868),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__53751),
            .ce(N__35458),
            .sr(N__53379));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_12_19_3  (
            .in0(N__35622),
            .in1(N__34861),
            .in2(_gnd_net_),
            .in3(N__34844),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__53751),
            .ce(N__35458),
            .sr(N__53379));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_12_19_4  (
            .in0(N__35588),
            .in1(N__34839),
            .in2(_gnd_net_),
            .in3(N__34820),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__53751),
            .ce(N__35458),
            .sr(N__53379));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_12_19_5  (
            .in0(N__35623),
            .in1(N__34813),
            .in2(_gnd_net_),
            .in3(N__34796),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__53751),
            .ce(N__35458),
            .sr(N__53379));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_12_19_6  (
            .in0(N__35589),
            .in1(N__34789),
            .in2(_gnd_net_),
            .in3(N__34772),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__53751),
            .ce(N__35458),
            .sr(N__53379));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_12_19_7  (
            .in0(N__35624),
            .in1(N__34765),
            .in2(_gnd_net_),
            .in3(N__34748),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__53751),
            .ce(N__35458),
            .sr(N__53379));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_12_20_0  (
            .in0(N__35602),
            .in1(N__34741),
            .in2(_gnd_net_),
            .in3(N__34724),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__53746),
            .ce(N__35475),
            .sr(N__53385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_12_20_1  (
            .in0(N__35618),
            .in1(N__34717),
            .in2(_gnd_net_),
            .in3(N__34700),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__53746),
            .ce(N__35475),
            .sr(N__53385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_12_20_2  (
            .in0(N__35599),
            .in1(N__34693),
            .in2(_gnd_net_),
            .in3(N__34676),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__53746),
            .ce(N__35475),
            .sr(N__53385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_12_20_3  (
            .in0(N__35615),
            .in1(N__35071),
            .in2(_gnd_net_),
            .in3(N__35054),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__53746),
            .ce(N__35475),
            .sr(N__53385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_12_20_4  (
            .in0(N__35600),
            .in1(N__35047),
            .in2(_gnd_net_),
            .in3(N__35030),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__53746),
            .ce(N__35475),
            .sr(N__53385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_12_20_5  (
            .in0(N__35616),
            .in1(N__35023),
            .in2(_gnd_net_),
            .in3(N__35006),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__53746),
            .ce(N__35475),
            .sr(N__53385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_12_20_6  (
            .in0(N__35601),
            .in1(N__34999),
            .in2(_gnd_net_),
            .in3(N__34982),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__53746),
            .ce(N__35475),
            .sr(N__53385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_12_20_7  (
            .in0(N__35617),
            .in1(N__34975),
            .in2(_gnd_net_),
            .in3(N__34958),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__53746),
            .ce(N__35475),
            .sr(N__53385));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_12_21_0  (
            .in0(N__35603),
            .in1(N__34951),
            .in2(_gnd_net_),
            .in3(N__34934),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__53741),
            .ce(N__35482),
            .sr(N__53391));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_12_21_1  (
            .in0(N__35611),
            .in1(N__34927),
            .in2(_gnd_net_),
            .in3(N__34910),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__53741),
            .ce(N__35482),
            .sr(N__53391));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_12_21_2  (
            .in0(N__35604),
            .in1(N__34903),
            .in2(_gnd_net_),
            .in3(N__34886),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__53741),
            .ce(N__35482),
            .sr(N__53391));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_12_21_3  (
            .in0(N__35612),
            .in1(N__35257),
            .in2(_gnd_net_),
            .in3(N__35240),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__53741),
            .ce(N__35482),
            .sr(N__53391));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_12_21_4  (
            .in0(N__35605),
            .in1(N__35233),
            .in2(_gnd_net_),
            .in3(N__35216),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__53741),
            .ce(N__35482),
            .sr(N__53391));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_12_21_5  (
            .in0(N__35613),
            .in1(N__35209),
            .in2(_gnd_net_),
            .in3(N__35192),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__53741),
            .ce(N__35482),
            .sr(N__53391));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_12_21_6  (
            .in0(N__35606),
            .in1(N__35185),
            .in2(_gnd_net_),
            .in3(N__35168),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__53741),
            .ce(N__35482),
            .sr(N__53391));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_12_21_7  (
            .in0(N__35614),
            .in1(N__35161),
            .in2(_gnd_net_),
            .in3(N__35144),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__53741),
            .ce(N__35482),
            .sr(N__53391));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_12_22_0  (
            .in0(N__35607),
            .in1(N__35137),
            .in2(_gnd_net_),
            .in3(N__35120),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__53736),
            .ce(N__35483),
            .sr(N__53401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_12_22_1  (
            .in0(N__35619),
            .in1(N__35113),
            .in2(_gnd_net_),
            .in3(N__35096),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__53736),
            .ce(N__35483),
            .sr(N__53401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_12_22_2  (
            .in0(N__35608),
            .in1(N__35093),
            .in2(_gnd_net_),
            .in3(N__35078),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__53736),
            .ce(N__35483),
            .sr(N__53401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_12_22_3  (
            .in0(N__35620),
            .in1(N__35662),
            .in2(_gnd_net_),
            .in3(N__35645),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__53736),
            .ce(N__35483),
            .sr(N__53401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_12_22_4  (
            .in0(N__35609),
            .in1(N__35641),
            .in2(_gnd_net_),
            .in3(N__35627),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__53736),
            .ce(N__35483),
            .sr(N__53401));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_22_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_12_22_5  (
            .in0(N__35495),
            .in1(N__35610),
            .in2(_gnd_net_),
            .in3(N__35498),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53736),
            .ce(N__35483),
            .sr(N__53401));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_12_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_12_23_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__35441),
            .in2(N__35420),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_12_23_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_12_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_12_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(N__35399),
            .in2(N__35381),
            .in3(N__35363),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_12_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_12_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__35360),
            .in2(N__35342),
            .in3(N__35324),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_12_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_12_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__35321),
            .in2(N__35303),
            .in3(N__35282),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_12_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_12_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__35279),
            .in2(N__35981),
            .in3(N__35264),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_12_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_12_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__35958),
            .in2(N__35849),
            .in3(N__35828),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_12_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_12_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__35825),
            .in2(N__35982),
            .in3(N__35810),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_12_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_12_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_12_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(N__35962),
            .in2(N__35807),
            .in3(N__35783),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_12_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_12_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__35963),
            .in2(N__35780),
            .in3(N__35762),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_12_24_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_12_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_12_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(N__35759),
            .in2(N__35983),
            .in3(N__35741),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_12_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_12_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(N__35738),
            .in2(N__35986),
            .in3(N__35723),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_12_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_12_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_12_24_3  (
            .in0(_gnd_net_),
            .in1(N__35720),
            .in2(N__35984),
            .in3(N__35705),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_12_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_12_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_12_24_4  (
            .in0(_gnd_net_),
            .in1(N__35702),
            .in2(N__35987),
            .in3(N__35687),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_12_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_12_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_12_24_5  (
            .in0(_gnd_net_),
            .in1(N__35684),
            .in2(N__35985),
            .in3(N__35669),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_12_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_12_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(N__35973),
            .in2(N__35900),
            .in3(N__35882),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_12_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_12_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_12_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35879),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_3.C_ON=1'b0;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53462),
            .lcout(GB_BUFFER_red_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_13_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_13_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_13_6_1  (
            .in0(N__35864),
            .in1(N__43781),
            .in2(_gnd_net_),
            .in3(N__40630),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(elapsed_time_ns_1_RNI24CN9_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_13_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_13_6_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35858),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_13_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_13_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_13_6_4  (
            .in0(N__40631),
            .in1(N__44213),
            .in2(_gnd_net_),
            .in3(N__37729),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37198),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_13_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_13_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37351),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_13_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_13_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__35855),
            .in2(N__37730),
            .in3(N__37483),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_13_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_13_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__36095),
            .in2(_gnd_net_),
            .in3(N__37471),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_13_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_13_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__37340),
            .in2(_gnd_net_),
            .in3(N__36089),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_13_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_13_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__38441),
            .in2(_gnd_net_),
            .in3(N__36074),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_13_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_13_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__36071),
            .in2(_gnd_net_),
            .in3(N__36053),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_13_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_13_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__37169),
            .in2(_gnd_net_),
            .in3(N__36038),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_13_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_13_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__37373),
            .in2(_gnd_net_),
            .in3(N__36023),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_13_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_13_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__37358),
            .in2(_gnd_net_),
            .in3(N__36008),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_13_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_13_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__37544),
            .in2(_gnd_net_),
            .in3(N__35990),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_13_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_13_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__37178),
            .in2(_gnd_net_),
            .in3(N__36227),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_13_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_13_8_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37394),
            .in3(N__36212),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_13_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_13_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__37421),
            .in2(_gnd_net_),
            .in3(N__36197),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_13_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_13_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__37490),
            .in2(_gnd_net_),
            .in3(N__36182),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_13_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_13_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__38366),
            .in2(_gnd_net_),
            .in3(N__36167),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_13_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_13_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__36164),
            .in2(_gnd_net_),
            .in3(N__36143),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_13_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_13_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__40493),
            .in2(_gnd_net_),
            .in3(N__36128),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_13_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_13_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__37565),
            .in2(_gnd_net_),
            .in3(N__36113),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_13_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_13_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__37559),
            .in2(_gnd_net_),
            .in3(N__36098),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_13_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_13_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__37415),
            .in2(_gnd_net_),
            .in3(N__36356),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_13_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_13_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__37427),
            .in2(_gnd_net_),
            .in3(N__36341),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_13_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_13_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__37508),
            .in2(_gnd_net_),
            .in3(N__36326),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_13_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_13_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__36323),
            .in2(_gnd_net_),
            .in3(N__36302),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_13_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_13_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__37529),
            .in2(_gnd_net_),
            .in3(N__36287),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_13_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_13_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__38492),
            .in2(_gnd_net_),
            .in3(N__36272),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_13_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_13_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__37553),
            .in2(_gnd_net_),
            .in3(N__36257),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_13_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_13_10_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37451),
            .in3(N__36242),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_13_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_13_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__38468),
            .in2(_gnd_net_),
            .in3(N__36545),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_13_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_13_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__37523),
            .in2(_gnd_net_),
            .in3(N__36530),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_13_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_13_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__37502),
            .in2(_gnd_net_),
            .in3(N__36515),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_13_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_13_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__36488),
            .in2(_gnd_net_),
            .in3(N__36500),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_13_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_13_10_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_13_10_6  (
            .in0(N__36497),
            .in1(N__37731),
            .in2(_gnd_net_),
            .in3(N__36491),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38429),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_28_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36478),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53790),
            .ce(N__37648),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_13_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_13_11_4 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_13_11_4  (
            .in0(N__36467),
            .in1(N__36434),
            .in2(_gnd_net_),
            .in3(N__36397),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_12_0 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_12_0  (
            .in0(N__39010),
            .in1(N__49750),
            .in2(N__39053),
            .in3(N__49948),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_12_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_13_12_1  (
            .in0(N__49946),
            .in1(N__38974),
            .in2(N__49766),
            .in3(N__38990),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_13_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_13_12_2 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_13_12_2  (
            .in0(N__38989),
            .in1(N__49944),
            .in2(N__38975),
            .in3(N__49746),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_13_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_13_12_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_13_12_3  (
            .in0(N__49945),
            .in1(N__39281),
            .in2(N__49765),
            .in3(N__39301),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_13_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_13_12_4 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_13_12_4  (
            .in0(N__38173),
            .in1(N__49751),
            .in2(N__38822),
            .in3(N__49950),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_12_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_13_12_5  (
            .in0(N__49947),
            .in1(N__38683),
            .in2(N__49767),
            .in3(N__38037),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_12_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_12_6  (
            .in0(N__38262),
            .in1(N__49752),
            .in2(N__38633),
            .in3(N__49949),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_13_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_13_12_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_13_12_7  (
            .in0(N__49951),
            .in1(N__38751),
            .in2(N__49768),
            .in3(N__38317),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_13_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_13_13_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_13_13_0  (
            .in0(N__49942),
            .in1(N__39349),
            .in2(N__49757),
            .in3(N__38193),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_13_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_13_13_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_13_13_1  (
            .in0(N__39350),
            .in1(N__49941),
            .in2(N__38195),
            .in3(N__49712),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39103),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53785),
            .ce(N__39076),
            .sr(N__53342));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_13_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_13_13_3 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_13_13_3  (
            .in0(N__38936),
            .in1(N__49713),
            .in2(N__38906),
            .in3(N__49940),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37821),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_13_5 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_13_5  (
            .in0(N__36590),
            .in1(_gnd_net_),
            .in2(N__36566),
            .in3(N__49936),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_13_6 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_13_6  (
            .in0(N__49714),
            .in1(N__38902),
            .in2(N__50021),
            .in3(N__38935),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_13_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_13_7  (
            .in0(N__36589),
            .in1(N__49935),
            .in2(_gnd_net_),
            .in3(N__36563),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38125),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36582),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_15_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_13_15_0  (
            .in0(N__49996),
            .in1(N__49553),
            .in2(N__38000),
            .in3(N__40735),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_13_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_13_15_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_13_15_1  (
            .in0(N__49554),
            .in1(N__49997),
            .in2(N__40739),
            .in3(N__37999),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_15_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_15_2  (
            .in0(N__49998),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49552),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_13_15_3  (
            .in0(N__39578),
            .in1(N__40734),
            .in2(_gnd_net_),
            .in3(N__37995),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_15_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_15_5  (
            .in0(N__39577),
            .in1(N__37822),
            .in2(_gnd_net_),
            .in3(N__36583),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39107),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53780),
            .ce(N__39075),
            .sr(N__53354));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45227),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53780),
            .ce(N__39075),
            .sr(N__53354));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_16_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_13_16_1  (
            .in0(N__49992),
            .in1(N__49717),
            .in2(N__38821),
            .in3(N__38174),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_16_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_13_16_2  (
            .in0(N__49719),
            .in1(N__49994),
            .in2(N__40804),
            .in3(N__38214),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38859),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_16_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_13_16_4  (
            .in0(N__49715),
            .in1(N__49995),
            .in2(N__39539),
            .in3(N__41273),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39419),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_6  (
            .in0(N__49718),
            .in1(N__49993),
            .in2(N__39725),
            .in3(N__39682),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_13_16_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_13_16_7  (
            .in0(N__49991),
            .in1(N__49716),
            .in2(N__38684),
            .in3(N__38039),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0  (
            .in0(N__49979),
            .in1(N__38146),
            .in2(N__45944),
            .in3(N__38124),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45191),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53770),
            .ce(N__39074),
            .sr(N__53365));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3  (
            .in0(N__38147),
            .in1(N__49978),
            .in2(N__38126),
            .in3(N__45943),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_13_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_13_17_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_13_17_6  (
            .in0(N__49980),
            .in1(N__49623),
            .in2(N__46427),
            .in3(N__38334),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_17_7 .LUT_INIT=16'b1111001111110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_17_7  (
            .in0(N__49622),
            .in1(N__49981),
            .in2(N__38341),
            .in3(N__46421),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_13_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_13_18_0 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_13_18_0  (
            .in0(N__39902),
            .in1(N__49727),
            .in2(N__39389),
            .in3(N__49986),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_2 .LUT_INIT=16'b1010000010101111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_18_2  (
            .in0(N__39458),
            .in1(N__49728),
            .in2(N__50141),
            .in3(N__39431),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_13_18_3  (
            .in0(N__49990),
            .in1(N__38866),
            .in2(N__49761),
            .in3(N__38242),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_18_4 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_13_18_4  (
            .in0(N__38867),
            .in1(N__49736),
            .in2(N__38243),
            .in3(N__49989),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_13_18_5  (
            .in0(N__49988),
            .in1(N__40805),
            .in2(N__49760),
            .in3(N__38219),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_13_18_6  (
            .in0(N__38318),
            .in1(N__49729),
            .in2(N__38759),
            .in3(N__49987),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_13_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_13_18_7  (
            .in0(N__49985),
            .in1(N__38625),
            .in2(N__49759),
            .in3(N__38270),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38533),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38287),
            .ce(),
            .sr(N__53380));
    defparam \pwm_generator_inst.un3_threshold_axb_8_LC_13_21_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_8_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_8_LC_13_21_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_8_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__36812),
            .in2(N__36791),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_13_21_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_13_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__36758),
            .in2(N__36740),
            .in3(N__36707),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_13_21_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_13_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__36704),
            .in2(N__36683),
            .in3(N__36650),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_13_21_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_13_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(N__36647),
            .in2(N__36629),
            .in3(N__36593),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_13_21_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_13_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(N__37163),
            .in2(N__36884),
            .in3(N__37130),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_13_21_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_13_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__36866),
            .in2(N__37127),
            .in3(N__37094),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_13_21_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_13_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(N__37091),
            .in2(N__36885),
            .in3(N__37064),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_13_21_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_13_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(N__36870),
            .in2(N__37061),
            .in3(N__37025),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_13_22_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_13_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__36886),
            .in2(N__37022),
            .in3(N__36989),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_13_22_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_13_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__36986),
            .in2(N__36897),
            .in3(N__36956),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_13_22_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_13_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__36953),
            .in2(N__36899),
            .in3(N__36920),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_13_22_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_13_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(N__36917),
            .in2(N__36898),
            .in3(N__37322),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_13_22_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_13_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37319),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_22_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_22_6  (
            .in0(N__53461),
            .in1(N__37300),
            .in2(_gnd_net_),
            .in3(N__37231),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37304),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53738),
            .ce(),
            .sr(N__53402));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_13_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_13_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_13_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40225),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53738),
            .ce(),
            .sr(N__53402));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_13_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_13_23_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_13_23_7  (
            .in0(N__40156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53738),
            .ce(),
            .sr(N__53402));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_14_5_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_14_5_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_14_5_0  (
            .in0(N__40605),
            .in1(N__37199),
            .in2(_gnd_net_),
            .in3(N__44000),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_14_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_14_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_14_5_1  (
            .in0(N__37187),
            .in1(N__43889),
            .in2(_gnd_net_),
            .in3(N__40604),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(elapsed_time_ns_1_RNITUBN9_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_14_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_14_5_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37181),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_14_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_14_6_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_14_6_0  (
            .in0(N__38386),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_6_1  (
            .in0(N__37403),
            .in1(N__43865),
            .in2(_gnd_net_),
            .in3(N__40582),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(elapsed_time_ns_1_RNIUVBN9_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_14_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_14_6_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37397),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_14_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_14_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_14_6_3  (
            .in0(N__43612),
            .in1(N__37382),
            .in2(_gnd_net_),
            .in3(N__40580),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_14_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_14_6_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37376),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_14_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_14_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_14_6_5  (
            .in0(N__37367),
            .in1(N__43583),
            .in2(_gnd_net_),
            .in3(N__40581),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(elapsed_time_ns_1_RNIK63T9_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_14_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_14_6_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37361),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_7  (
            .in0(N__37352),
            .in1(N__40583),
            .in2(_gnd_net_),
            .in3(N__43655),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_14_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_14_7_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_14_7_0  (
            .in0(N__38398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_14_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_14_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_14_7_1  (
            .in0(N__38581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_14_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_14_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_14_7_2  (
            .in0(N__37484),
            .in1(N__40409),
            .in2(_gnd_net_),
            .in3(N__40619),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_14_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_14_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_14_7_3  (
            .in0(N__40620),
            .in1(N__37472),
            .in2(_gnd_net_),
            .in3(N__40391),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_14_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_14_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_14_7_4  (
            .in0(N__37439),
            .in1(N__44042),
            .in2(_gnd_net_),
            .in3(N__40621),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_14_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_14_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_14_7_6  (
            .in0(N__37460),
            .in1(N__43910),
            .in2(_gnd_net_),
            .in3(N__40618),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(elapsed_time_ns_1_RNI47DN9_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_14_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_14_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37454),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_14_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_14_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37438),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_14_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_14_8_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_14_8_1  (
            .in0(N__38353),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_14_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_14_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_14_8_2  (
            .in0(N__38569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_14_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_14_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_14_8_3  (
            .in0(N__40622),
            .in1(N__37409),
            .in2(_gnd_net_),
            .in3(N__43556),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(elapsed_time_ns_1_RNIL73T9_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_14_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_14_8_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37547),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_14_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_14_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_14_8_6  (
            .in0(N__37538),
            .in1(N__43979),
            .in2(_gnd_net_),
            .in3(N__40623),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(elapsed_time_ns_1_RNI14DN9_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_14_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_14_8_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37532),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_14_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_14_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38455),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_14_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_14_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_14_9_2  (
            .in0(N__40625),
            .in1(N__37517),
            .in2(_gnd_net_),
            .in3(N__44021),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(elapsed_time_ns_1_RNIV1DN9_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_14_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_14_9_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37511),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_14_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_14_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40649),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_14_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_14_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_14_9_5  (
            .in0(N__37496),
            .in1(N__43742),
            .in2(_gnd_net_),
            .in3(N__40624),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(elapsed_time_ns_1_RNI46CN9_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_14_9_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37568),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_14_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_14_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38512),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_14_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_14_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38704),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38604),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38952),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38655),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39032),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38730),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41696),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39263),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42828),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_14_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_14_11_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_14_11_4  (
            .in0(N__50059),
            .in1(N__40851),
            .in2(N__49769),
            .in3(N__38092),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49785),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_14_11_6  (
            .in0(N__39738),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_11_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__38922),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_14_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_14_12_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_0_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__37736),
            .in2(_gnd_net_),
            .in3(N__37685),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53791),
            .ce(N__37643),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41801),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_12_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__38790),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39190),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39363),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39495),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39699),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39129),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__37829),
            .in2(N__37823),
            .in3(N__37820),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__37796),
            .in2(_gnd_net_),
            .in3(N__37787),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__37784),
            .in2(_gnd_net_),
            .in3(N__37775),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__37772),
            .in2(_gnd_net_),
            .in3(N__37763),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__37760),
            .in2(_gnd_net_),
            .in3(N__37751),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__37748),
            .in2(_gnd_net_),
            .in3(N__37739),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__37919),
            .in2(_gnd_net_),
            .in3(N__37910),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__37907),
            .in2(_gnd_net_),
            .in3(N__37898),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__39317),
            .in2(_gnd_net_),
            .in3(N__37895),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__37892),
            .in2(_gnd_net_),
            .in3(N__37883),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__37880),
            .in2(_gnd_net_),
            .in3(N__37871),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__37868),
            .in2(_gnd_net_),
            .in3(N__37859),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__37856),
            .in2(_gnd_net_),
            .in3(N__37844),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__37841),
            .in2(_gnd_net_),
            .in3(N__37832),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__40829),
            .in2(_gnd_net_),
            .in3(N__38018),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__38015),
            .in2(_gnd_net_),
            .in3(N__38006),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__40751),
            .in2(_gnd_net_),
            .in3(N__38003),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__40709),
            .in2(_gnd_net_),
            .in3(N__37985),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__37982),
            .in2(_gnd_net_),
            .in3(N__37970),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__37967),
            .in2(_gnd_net_),
            .in3(N__37958),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__37955),
            .in2(_gnd_net_),
            .in3(N__37946),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__37943),
            .in2(_gnd_net_),
            .in3(N__37934),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__37931),
            .in2(_gnd_net_),
            .in3(N__37922),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__40817),
            .in2(_gnd_net_),
            .in3(N__38072),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__40763),
            .in2(_gnd_net_),
            .in3(N__38069),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__38066),
            .in2(_gnd_net_),
            .in3(N__38060),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__40697),
            .in2(_gnd_net_),
            .in3(N__38057),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__41237),
            .in2(_gnd_net_),
            .in3(N__38054),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__38051),
            .in2(_gnd_net_),
            .in3(N__38045),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38042),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_14_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_14_16_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_14_16_6  (
            .in0(N__49639),
            .in1(N__50049),
            .in2(N__38096),
            .in3(N__40861),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_16_7  (
            .in0(N__39585),
            .in1(N__38673),
            .in2(_gnd_net_),
            .in3(N__38038),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_17_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_17_0  (
            .in0(N__39481),
            .in1(N__50096),
            .in2(N__49758),
            .in3(N__39515),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_17_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_14_17_1  (
            .in0(N__50095),
            .in1(N__49723),
            .in2(N__39218),
            .in3(N__39241),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_17_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_17_2  (
            .in0(N__39348),
            .in1(N__39653),
            .in2(_gnd_net_),
            .in3(N__38194),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_14_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_14_17_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_14_17_3  (
            .in0(N__39657),
            .in1(_gnd_net_),
            .in2(N__41722),
            .in3(N__41745),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_17_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_17_4  (
            .in0(N__38808),
            .in1(N__39655),
            .in2(_gnd_net_),
            .in3(N__38172),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_17_5  (
            .in0(N__39656),
            .in1(N__39754),
            .in2(_gnd_net_),
            .in3(N__39778),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_14_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_14_17_6 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_14_17_6  (
            .in0(N__38140),
            .in1(N__38120),
            .in2(_gnd_net_),
            .in3(N__39652),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_17_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_17_7  (
            .in0(N__39654),
            .in1(_gnd_net_),
            .in2(N__42850),
            .in3(N__42876),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_14_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_14_18_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_14_18_0  (
            .in0(N__39635),
            .in1(_gnd_net_),
            .in2(N__40862),
            .in3(N__38091),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_14_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_14_18_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_14_18_1  (
            .in0(N__39214),
            .in1(N__39637),
            .in2(_gnd_net_),
            .in3(N__39240),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_14_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_14_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_14_18_2  (
            .in0(N__39633),
            .in1(N__38629),
            .in2(_gnd_net_),
            .in3(N__38269),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_14_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_14_18_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_14_18_3  (
            .in0(N__41820),
            .in1(N__39636),
            .in2(_gnd_net_),
            .in3(N__41776),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_14_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_14_18_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_14_18_4  (
            .in0(N__39639),
            .in1(N__39174),
            .in2(_gnd_net_),
            .in3(N__39147),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_18_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_18_5  (
            .in0(N__39381),
            .in1(N__39634),
            .in2(_gnd_net_),
            .in3(N__39901),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_14_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_14_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_14_18_6  (
            .in0(N__39638),
            .in1(N__39513),
            .in2(_gnd_net_),
            .in3(N__39480),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_14_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_14_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_14_19_0  (
            .in0(N__50118),
            .in1(N__38865),
            .in2(_gnd_net_),
            .in3(N__38238),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_14_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_14_19_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_14_19_1  (
            .in0(N__42987),
            .in1(N__39664),
            .in2(_gnd_net_),
            .in3(N__42943),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_19_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_19_2  (
            .in0(N__50117),
            .in1(N__40797),
            .in2(_gnd_net_),
            .in3(N__38215),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_14_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_14_19_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_14_19_3  (
            .in0(N__39430),
            .in1(N__50121),
            .in2(_gnd_net_),
            .in3(N__39451),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4 .LUT_INIT=16'b1100010111000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_19_4  (
            .in0(N__39148),
            .in1(N__39179),
            .in2(N__50135),
            .in3(N__49624),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_19_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_14_19_5  (
            .in0(N__41272),
            .in1(N__50120),
            .in2(_gnd_net_),
            .in3(N__39538),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_14_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_14_19_6 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_14_19_6  (
            .in0(N__41674),
            .in1(_gnd_net_),
            .in2(N__39665),
            .in3(N__41634),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_19_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__50119),
            .in2(N__43066),
            .in3(N__43107),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_14_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_14_20_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__50091),
            .in2(_gnd_net_),
            .in3(N__38342),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_20_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_14_20_4  (
            .in0(N__38310),
            .in1(N__39660),
            .in2(_gnd_net_),
            .in3(N__38752),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_14_21_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_14_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_14_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38532),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38288),
            .ce(),
            .sr(N__53381));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_5_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_5_2  (
            .in0(N__43582),
            .in1(N__40421),
            .in2(N__43613),
            .in3(N__40415),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_15_6_1  (
            .in0(N__43676),
            .in1(N__38276),
            .in2(_gnd_net_),
            .in3(N__40577),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(elapsed_time_ns_1_RNIG23T9_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_15_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_15_6_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38444),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_15_6_3  (
            .in0(N__44234),
            .in1(N__38425),
            .in2(_gnd_net_),
            .in3(N__40579),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_15_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_15_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_15_6_4  (
            .in0(N__40679),
            .in1(N__40664),
            .in2(N__40658),
            .in3(N__40685),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_6_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_6_5  (
            .in0(N__44209),
            .in1(N__40670),
            .in2(N__38411),
            .in3(N__38408),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_6_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_6_6  (
            .in0(N__38399),
            .in1(_gnd_net_),
            .in2(N__38402),
            .in3(N__43694),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_6_7  (
            .in0(N__38387),
            .in1(N__43634),
            .in2(_gnd_net_),
            .in3(N__40578),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0  (
            .in0(N__43802),
            .in1(N__38375),
            .in2(_gnd_net_),
            .in3(N__40606),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(elapsed_time_ns_1_RNI13CN9_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_15_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_15_7_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38369),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_15_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_15_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_15_7_3  (
            .in0(N__40607),
            .in1(N__38354),
            .in2(_gnd_net_),
            .in3(N__43844),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_15_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_15_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_15_7_5  (
            .in0(N__40610),
            .in1(N__38480),
            .in2(_gnd_net_),
            .in3(N__44291),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_15_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_15_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_15_7_6  (
            .in0(N__38582),
            .in1(N__43823),
            .in2(_gnd_net_),
            .in3(N__40608),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_7_7  (
            .in0(N__40609),
            .in1(N__38570),
            .in2(_gnd_net_),
            .in3(N__44063),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_8_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_8_0  (
            .in0(N__41105),
            .in1(N__38551),
            .in2(_gnd_net_),
            .in3(N__41141),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_8_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_8_1  (
            .in0(N__40627),
            .in1(N__38513),
            .in2(_gnd_net_),
            .in3(N__43718),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_8_2  (
            .in0(N__38501),
            .in1(N__43955),
            .in2(_gnd_net_),
            .in3(N__40626),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(elapsed_time_ns_1_RNI25DN9_0_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_15_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_15_8_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38495),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_15_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38479),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_15_9_1  (
            .in0(N__40629),
            .in1(N__38456),
            .in2(_gnd_net_),
            .in3(N__44270),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_15_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_15_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_15_9_4  (
            .in0(N__38705),
            .in1(N__43934),
            .in2(_gnd_net_),
            .in3(N__40628),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__45151),
            .in2(N__45223),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__53814),
            .ce(N__39080),
            .sr(N__53327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__45127),
            .in2(N__45190),
            .in3(N__38693),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__53814),
            .ce(N__39080),
            .sr(N__53327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__45152),
            .in2(N__45103),
            .in3(N__38690),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__53814),
            .ce(N__39080),
            .sr(N__53327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__45128),
            .in2(N__45073),
            .in3(N__38687),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__53814),
            .ce(N__39080),
            .sr(N__53327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__45040),
            .in2(N__45104),
            .in3(N__38639),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__53814),
            .ce(N__39080),
            .sr(N__53327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__45643),
            .in2(N__45074),
            .in3(N__38636),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__53814),
            .ce(N__39080),
            .sr(N__53327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__45616),
            .in2(N__45044),
            .in3(N__38588),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__53814),
            .ce(N__39080),
            .sr(N__53327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__45644),
            .in2(N__45583),
            .in3(N__38585),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__53814),
            .ce(N__39080),
            .sr(N__53327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__45541),
            .in2(N__45620),
            .in3(N__38825),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__53805),
            .ce(N__39079),
            .sr(N__53329));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__45514),
            .in2(N__45584),
            .in3(N__38774),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__53805),
            .ce(N__39079),
            .sr(N__53329));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__45490),
            .in2(N__45545),
            .in3(N__38771),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__53805),
            .ce(N__39079),
            .sr(N__53329));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__45515),
            .in2(N__45466),
            .in3(N__38768),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__53805),
            .ce(N__39079),
            .sr(N__53329));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__45491),
            .in2(N__45436),
            .in3(N__38765),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__53805),
            .ce(N__39079),
            .sr(N__53329));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__45910),
            .in2(N__45467),
            .in3(N__38762),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__53805),
            .ce(N__39079),
            .sr(N__53329));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__45883),
            .in2(N__45437),
            .in3(N__38714),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__53805),
            .ce(N__39079),
            .sr(N__53329));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__45911),
            .in2(N__45850),
            .in3(N__38711),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__53805),
            .ce(N__39079),
            .sr(N__53329));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__45808),
            .in2(N__45887),
            .in3(N__38708),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__53799),
            .ce(N__39078),
            .sr(N__53335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__45781),
            .in2(N__45851),
            .in3(N__38888),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__53799),
            .ce(N__39078),
            .sr(N__53335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__45754),
            .in2(N__45812),
            .in3(N__38885),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__53799),
            .ce(N__39078),
            .sr(N__53335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__45782),
            .in2(N__45727),
            .in3(N__38882),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__53799),
            .ce(N__39078),
            .sr(N__53335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__45694),
            .in2(N__45758),
            .in3(N__38879),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__53799),
            .ce(N__39078),
            .sr(N__53335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__45667),
            .in2(N__45728),
            .in3(N__38876),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__53799),
            .ce(N__39078),
            .sr(N__53335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__46165),
            .in2(N__45698),
            .in3(N__38873),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__53799),
            .ce(N__39078),
            .sr(N__53335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__45668),
            .in2(N__46132),
            .in3(N__38870),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__53799),
            .ce(N__39078),
            .sr(N__53335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__46093),
            .in2(N__46169),
            .in3(N__38831),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__53792),
            .ce(N__39077),
            .sr(N__53337));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__46069),
            .in2(N__46133),
            .in3(N__38828),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__53792),
            .ce(N__39077),
            .sr(N__53337));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__46094),
            .in2(N__46046),
            .in3(N__39116),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__53792),
            .ce(N__39077),
            .sr(N__53337));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__46070),
            .in2(N__46016),
            .in3(N__39113),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__53792),
            .ce(N__39077),
            .sr(N__53337));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39110),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39096),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53792),
            .ce(N__39077),
            .sr(N__53337));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_14_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_14_0  (
            .in0(N__39280),
            .in1(N__39649),
            .in2(_gnd_net_),
            .in3(N__39297),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_14_1  (
            .in0(N__39651),
            .in1(N__39042),
            .in2(_gnd_net_),
            .in3(N__39006),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_14_2 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_14_2  (
            .in0(N__38988),
            .in1(N__39650),
            .in2(_gnd_net_),
            .in3(N__38965),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_14_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_14_3  (
            .in0(N__39648),
            .in1(N__38929),
            .in2(_gnd_net_),
            .in3(N__38901),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_14_4 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_15_14_4  (
            .in0(N__49649),
            .in1(N__39777),
            .in2(N__50126),
            .in3(N__39753),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_14_5 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_14_5  (
            .in0(N__41749),
            .in1(N__50111),
            .in2(N__41723),
            .in3(N__49650),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39339),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_15_14_7  (
            .in0(N__39311),
            .in1(_gnd_net_),
            .in2(N__42703),
            .in3(N__39872),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_15_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_15_0  (
            .in0(N__49558),
            .in1(N__50089),
            .in2(N__39724),
            .in3(N__39683),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_15_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_15_15_1  (
            .in0(N__50087),
            .in1(N__49559),
            .in2(N__41821),
            .in3(N__41775),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_15_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_15_15_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_15_15_2  (
            .in0(N__49555),
            .in1(N__50083),
            .in2(N__39305),
            .in3(N__39279),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_15_3 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_15_15_3  (
            .in0(N__50086),
            .in1(N__41670),
            .in2(N__41638),
            .in3(N__49563),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_15_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_15_15_4  (
            .in0(N__49561),
            .in1(N__50088),
            .in2(N__39242),
            .in3(N__39213),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_15_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_15_5  (
            .in0(N__50090),
            .in1(N__49560),
            .in2(N__39178),
            .in3(N__39149),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_15_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_15_15_6  (
            .in0(N__49557),
            .in1(N__50085),
            .in2(N__39779),
            .in3(N__39755),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_15_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_15_7  (
            .in0(N__50084),
            .in1(N__49556),
            .in2(N__42880),
            .in3(N__42843),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_16_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_16_0  (
            .in0(N__39658),
            .in1(N__49792),
            .in2(_gnd_net_),
            .in3(N__50158),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_16_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_16_1  (
            .in0(N__39708),
            .in1(N__39681),
            .in2(_gnd_net_),
            .in3(N__39659),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_16_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_16_2  (
            .in0(N__42991),
            .in1(N__50099),
            .in2(N__49708),
            .in3(N__42942),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_16_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_15_16_3  (
            .in0(N__50101),
            .in1(N__41268),
            .in2(N__49706),
            .in3(N__39537),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_16_4 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_15_16_4  (
            .in0(N__39514),
            .in1(N__50098),
            .in2(N__39482),
            .in3(N__49634),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_16_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_16_5  (
            .in0(N__50100),
            .in1(N__43108),
            .in2(N__49705),
            .in3(N__43059),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_16_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_16_6  (
            .in0(N__39450),
            .in1(N__49635),
            .in2(N__39429),
            .in3(N__50102),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_16_7  (
            .in0(N__50097),
            .in1(N__39385),
            .in2(N__49707),
            .in3(N__39897),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__39871),
            .in2(N__46419),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__42416),
            .in2(N__39848),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__39836),
            .in2(N__42549),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__42420),
            .in2(N__39827),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__39818),
            .in2(N__42550),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__42424),
            .in2(N__39809),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__39797),
            .in2(N__42551),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__42428),
            .in2(N__39791),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__42542),
            .in2(N__39962),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__39953),
            .in2(N__42623),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__42530),
            .in2(N__39947),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__39938),
            .in2(N__42620),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__42534),
            .in2(N__39932),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__39923),
            .in2(N__42621),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__42538),
            .in2(N__39917),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__39908),
            .in2(N__42622),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__42514),
            .in2(N__40049),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__40037),
            .in2(N__42616),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__42518),
            .in2(N__40031),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__40013),
            .in2(N__42617),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__42522),
            .in2(N__40007),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__39998),
            .in2(N__42618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__42526),
            .in2(N__39992),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__39977),
            .in2(N__42619),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__42501),
            .in2(N__39971),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__40103),
            .in2(N__42613),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__42505),
            .in2(N__40097),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__40088),
            .in2(N__42614),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__42509),
            .in2(N__40082),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(N__40073),
            .in2(N__42615),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__42513),
            .in2(N__40067),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(N__50125),
            .in2(_gnd_net_),
            .in3(N__40058),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_15_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_15_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__40055),
            .in2(_gnd_net_),
            .in3(N__46805),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_15_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_15_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__47159),
            .in2(_gnd_net_),
            .in3(N__40130),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__53759),
            .ce(),
            .sr(N__53374));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_15_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_15_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__47138),
            .in2(_gnd_net_),
            .in3(N__40127),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__53759),
            .ce(),
            .sr(N__53374));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_15_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_15_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__47117),
            .in2(_gnd_net_),
            .in3(N__40124),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__53759),
            .ce(),
            .sr(N__53374));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_15_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_15_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_15_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__47096),
            .in2(_gnd_net_),
            .in3(N__40121),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__53759),
            .ce(),
            .sr(N__53374));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_15_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_15_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_15_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__47075),
            .in2(_gnd_net_),
            .in3(N__40118),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__53759),
            .ce(),
            .sr(N__53374));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_15_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_15_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_15_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__47054),
            .in2(_gnd_net_),
            .in3(N__40115),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__53759),
            .ce(),
            .sr(N__53374));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_15_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_15_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__47033),
            .in2(_gnd_net_),
            .in3(N__40112),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__53759),
            .ce(),
            .sr(N__53374));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_15_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_15_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__47012),
            .in2(_gnd_net_),
            .in3(N__40109),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__53753),
            .ce(),
            .sr(N__53382));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_15_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_15_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_15_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__47339),
            .in2(_gnd_net_),
            .in3(N__40106),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__53753),
            .ce(),
            .sr(N__53382));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_15_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_15_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__47318),
            .in2(_gnd_net_),
            .in3(N__40181),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__53753),
            .ce(),
            .sr(N__53382));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_15_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_15_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__47297),
            .in2(_gnd_net_),
            .in3(N__40178),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__53753),
            .ce(),
            .sr(N__53382));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_15_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_15_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__47273),
            .in2(_gnd_net_),
            .in3(N__40175),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__53753),
            .ce(),
            .sr(N__53382));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_15_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_15_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__47249),
            .in2(_gnd_net_),
            .in3(N__40172),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__53753),
            .ce(),
            .sr(N__53382));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_15_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_15_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__47225),
            .in2(_gnd_net_),
            .in3(N__40169),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__53753),
            .ce(),
            .sr(N__53382));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_15_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_15_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(N__47204),
            .in2(_gnd_net_),
            .in3(N__40166),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__53753),
            .ce(),
            .sr(N__53382));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_15_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_15_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_15_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__47180),
            .in2(_gnd_net_),
            .in3(N__40163),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__53748),
            .ce(),
            .sr(N__53386));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_15_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_15_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__47513),
            .in2(_gnd_net_),
            .in3(N__40136),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__53748),
            .ce(),
            .sr(N__53386));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_15_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_15_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_15_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__47486),
            .in2(_gnd_net_),
            .in3(N__40133),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__53748),
            .ce(),
            .sr(N__53386));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_15_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_15_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__47459),
            .in2(_gnd_net_),
            .in3(N__40208),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__53748),
            .ce(),
            .sr(N__53386));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_15_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_15_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_15_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__47438),
            .in2(_gnd_net_),
            .in3(N__40205),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__53748),
            .ce(),
            .sr(N__53386));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_15_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_15_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_15_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__47417),
            .in2(_gnd_net_),
            .in3(N__40202),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__53748),
            .ce(),
            .sr(N__53386));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_15_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_15_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_15_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__47393),
            .in2(_gnd_net_),
            .in3(N__40199),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__53748),
            .ce(),
            .sr(N__53386));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_15_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_15_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_15_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__47372),
            .in2(_gnd_net_),
            .in3(N__40196),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__53748),
            .ce(),
            .sr(N__53386));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_15_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_15_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_15_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__47831),
            .in2(_gnd_net_),
            .in3(N__40193),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__53743),
            .ce(),
            .sr(N__53392));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_15_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_15_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_15_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__47810),
            .in2(_gnd_net_),
            .in3(N__40190),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__53743),
            .ce(),
            .sr(N__53392));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_15_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_15_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__47783),
            .in2(_gnd_net_),
            .in3(N__40187),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .clk(N__53743),
            .ce(),
            .sr(N__53392));
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_15_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_15_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_15_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_27_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__47762),
            .in2(_gnd_net_),
            .in3(N__40184),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .clk(N__53743),
            .ce(),
            .sr(N__53392));
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_15_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_15_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_15_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_28_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__47738),
            .in2(_gnd_net_),
            .in3(N__40370),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .clk(N__53743),
            .ce(),
            .sr(N__53392));
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_15_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_15_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_15_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_29_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__47723),
            .in2(_gnd_net_),
            .in3(N__40367),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .clk(N__53743),
            .ce(),
            .sr(N__53392));
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_15_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_15_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_15_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_30_LC_15_24_6  (
            .in0(_gnd_net_),
            .in1(N__43397),
            .in2(_gnd_net_),
            .in3(N__40364),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ),
            .clk(N__53743),
            .ce(),
            .sr(N__53392));
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_15_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_15_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_15_24_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_31_LC_15_24_7  (
            .in0(_gnd_net_),
            .in1(N__47705),
            .in2(_gnd_net_),
            .in3(N__40361),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53743),
            .ce(),
            .sr(N__53392));
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_15_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_15_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_15_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_30_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40351),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53739),
            .ce(),
            .sr(N__53403));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_15_25_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_15_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_15_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40327),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53739),
            .ce(),
            .sr(N__53403));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_15_25_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_15_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_15_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40300),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53739),
            .ce(),
            .sr(N__53403));
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_15_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_15_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_15_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_29_LC_15_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40273),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53739),
            .ce(),
            .sr(N__53403));
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_15_26_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_15_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_15_26_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_27_LC_15_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40255),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53732),
            .ce(),
            .sr(N__53407));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_15_26_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_15_26_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_15_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40474),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53732),
            .ce(),
            .sr(N__53407));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_15_26_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_15_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_15_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40450),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53732),
            .ce(),
            .sr(N__53407));
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_15_26_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_15_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_15_26_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_31_LC_15_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40430),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53732),
            .ce(),
            .sr(N__53407));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_15_27_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_15_27_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_15_27_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_15_27_2  (
            .in0(N__52423),
            .in1(N__48188),
            .in2(_gnd_net_),
            .in3(N__52240),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53730),
            .ce(),
            .sr(N__53411));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_28_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_28_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_28_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_15_28_4  (
            .in0(N__52417),
            .in1(N__52196),
            .in2(_gnd_net_),
            .in3(N__48350),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53728),
            .ce(),
            .sr(N__53414));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_15_28_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_15_28_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_15_28_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_15_28_6  (
            .in0(N__52416),
            .in1(N__48134),
            .in2(_gnd_net_),
            .in3(N__52197),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53728),
            .ce(),
            .sr(N__53414));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_16_4_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_16_4_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_16_4_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_16_4_0  (
            .in0(N__43687),
            .in1(N__43669),
            .in2(N__40387),
            .in3(N__40402),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_4_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_4_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_4_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_4_2  (
            .in0(N__43627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43648),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_16_4_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_16_4_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_16_4_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_16_4_3  (
            .in0(N__44150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53852),
            .ce(N__44192),
            .sr(N__53314));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_4_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_4_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_4_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_4_5  (
            .in0(N__44119),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53852),
            .ce(N__44192),
            .sr(N__53314));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_5_2  (
            .in0(N__43774),
            .in1(N__43732),
            .in2(N__43714),
            .in3(N__43756),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_5_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_5_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_5_4  (
            .in0(N__44014),
            .in1(N__44035),
            .in2(N__43999),
            .in3(N__44056),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_16_5_5  (
            .in0(N__43885),
            .in1(N__43858),
            .in2(N__43552),
            .in3(N__43837),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_5_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_5_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_5_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_16_5_6  (
            .in0(_gnd_net_),
            .in1(N__43795),
            .in2(N__40673),
            .in3(N__43816),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_6_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_6_1  (
            .in0(N__44248),
            .in1(N__43948),
            .in2(N__43975),
            .in3(N__44230),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_16_6_5  (
            .in0(N__44284),
            .in1(N__43903),
            .in2(N__43930),
            .in3(N__44263),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_16_7_4  (
            .in0(N__40617),
            .in1(N__40645),
            .in2(_gnd_net_),
            .in3(N__44249),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_7_5  (
            .in0(N__40502),
            .in1(N__43760),
            .in2(_gnd_net_),
            .in3(N__40616),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(elapsed_time_ns_1_RNI35CN9_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_7_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40496),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__41104),
            .in2(_gnd_net_),
            .in3(N__41140),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_165_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41103),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_16_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_16_12_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_16_12_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_0_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__41078),
            .in2(_gnd_net_),
            .in3(N__41021),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53806),
            .ce(N__40967),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40845),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42968),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40779),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41657),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_12_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__40720),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43088),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41255),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__42796),
            .in2(N__45983),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__45931),
            .in2(N__41225),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__49487),
            .in2(N__41207),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_16_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_16_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__49157),
            .in2(N__49612),
            .in3(N__41195),
            .lcout(\current_shift_inst.un38_control_input_0_s1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_16_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_16_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__49491),
            .in2(N__41192),
            .in3(N__41180),
            .lcout(\current_shift_inst.un38_control_input_0_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_16_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_16_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__41177),
            .in2(N__49613),
            .in3(N__41165),
            .lcout(\current_shift_inst.un38_control_input_0_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_16_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_16_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__49495),
            .in2(N__41162),
            .in3(N__41144),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_16_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_16_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(N__41393),
            .in2(N__49614),
            .in3(N__41384),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_16_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_16_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__49326),
            .in2(N__41381),
            .in3(N__41363),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_16_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_16_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__41360),
            .in2(N__49502),
            .in3(N__41348),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_16_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_16_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__49330),
            .in2(N__42812),
            .in3(N__41345),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_16_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_16_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__41342),
            .in2(N__49503),
            .in3(N__41330),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_16_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_16_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__49334),
            .in2(N__41327),
            .in3(N__41312),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_16_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_16_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__41309),
            .in2(N__49504),
            .in3(N__41303),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_16_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_16_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__49338),
            .in2(N__41300),
            .in3(N__41291),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_16_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_16_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(N__41288),
            .in2(N__49505),
            .in3(N__41276),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_16_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_16_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__49404),
            .in2(N__41486),
            .in3(N__41471),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_16_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_16_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__41468),
            .in2(N__49545),
            .in3(N__41462),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_16_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_16_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__49408),
            .in2(N__41459),
            .in3(N__41447),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_16_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_16_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__41444),
            .in2(N__49546),
            .in3(N__41438),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__49412),
            .in2(N__41435),
            .in3(N__41426),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__41423),
            .in2(N__49547),
            .in3(N__41417),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__49416),
            .in2(N__41414),
            .in3(N__41405),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__41402),
            .in2(N__49548),
            .in3(N__41396),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__49420),
            .in2(N__41591),
            .in3(N__41582),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__41579),
            .in2(N__49549),
            .in3(N__41567),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__49424),
            .in2(N__41564),
            .in3(N__41549),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__41546),
            .in2(N__49550),
            .in3(N__41540),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__49428),
            .in2(N__41537),
            .in3(N__41528),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(N__41525),
            .in2(N__49551),
            .in3(N__41519),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_16_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_16_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(N__49432),
            .in2(N__41516),
            .in3(N__41501),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_16_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_16_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_16_16_7  (
            .in0(N__49433),
            .in1(N__50103),
            .in2(_gnd_net_),
            .in3(N__41498),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_17_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_17_0  (
            .in0(N__41495),
            .in1(N__46706),
            .in2(_gnd_net_),
            .in3(N__47680),
            .lcout(\current_shift_inst.control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_17_1 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_17_1  (
            .in0(N__50104),
            .in1(N__49539),
            .in2(N__42887),
            .in3(N__42851),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_17_3  (
            .in0(N__42800),
            .in1(N__42552),
            .in2(_gnd_net_),
            .in3(N__46420),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_16_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_16_17_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_16_17_4  (
            .in0(N__41831),
            .in1(N__46898),
            .in2(_gnd_net_),
            .in3(N__47681),
            .lcout(\current_shift_inst.control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_5  (
            .in0(N__50107),
            .in1(N__49540),
            .in2(N__41825),
            .in3(N__41780),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_16_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_16_17_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_16_17_6  (
            .in0(N__49541),
            .in1(N__50105),
            .in2(N__41753),
            .in3(N__41718),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_16_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_16_17_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_16_17_7  (
            .in0(N__50106),
            .in1(N__49542),
            .in2(N__41678),
            .in3(N__41639),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_18_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_18_0  (
            .in0(N__47663),
            .in1(N__41609),
            .in2(_gnd_net_),
            .in3(N__46943),
            .lcout(\current_shift_inst.control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_18_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_18_1  (
            .in0(N__47671),
            .in1(N__41600),
            .in2(_gnd_net_),
            .in3(N__46682),
            .lcout(\current_shift_inst.control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_18_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_18_2  (
            .in0(N__49543),
            .in1(N__50137),
            .in2(N__43115),
            .in3(N__43067),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_16_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_16_18_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_16_18_3  (
            .in0(N__46754),
            .in1(N__43037),
            .in2(_gnd_net_),
            .in3(N__47662),
            .lcout(\current_shift_inst.control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_18_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_18_4  (
            .in0(N__47661),
            .in1(N__46433),
            .in2(_gnd_net_),
            .in3(N__43028),
            .lcout(\current_shift_inst.control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_18_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_18_5  (
            .in0(N__46478),
            .in1(N__43016),
            .in2(_gnd_net_),
            .in3(N__47659),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_16_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_16_18_6 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_16_18_6  (
            .in0(N__47660),
            .in1(_gnd_net_),
            .in2(N__43007),
            .in3(N__46448),
            .lcout(\current_shift_inst.control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_18_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_18_7  (
            .in0(N__50136),
            .in1(N__49544),
            .in2(N__42992),
            .in3(N__42947),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_16_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_16_19_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_16_19_0  (
            .in0(N__42920),
            .in1(N__46328),
            .in2(_gnd_net_),
            .in3(N__47617),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_16_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_16_19_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_16_19_1  (
            .in0(N__47618),
            .in1(N__46301),
            .in2(_gnd_net_),
            .in3(N__42908),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_16_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_16_19_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_16_19_2  (
            .in0(N__42896),
            .in1(N__46271),
            .in2(_gnd_net_),
            .in3(N__47619),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_16_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_16_19_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_16_19_3  (
            .in0(N__47620),
            .in1(N__46244),
            .in2(_gnd_net_),
            .in3(N__43187),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_19_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_19_4  (
            .in0(N__43178),
            .in1(N__46985),
            .in2(_gnd_net_),
            .in3(N__47624),
            .lcout(\current_shift_inst.control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_16_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_16_19_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_16_19_5  (
            .in0(N__47623),
            .in1(N__43166),
            .in2(_gnd_net_),
            .in3(N__46604),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_16_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_16_19_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_16_19_6  (
            .in0(N__43157),
            .in1(N__46184),
            .in2(_gnd_net_),
            .in3(N__47622),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_16_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_16_19_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_16_19_7  (
            .in0(N__47621),
            .in1(N__46211),
            .in2(_gnd_net_),
            .in3(N__43148),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_20_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_20_0  (
            .in0(N__47614),
            .in1(N__43139),
            .in2(_gnd_net_),
            .in3(N__46556),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_20_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_20_1  (
            .in0(N__43127),
            .in1(N__46358),
            .in2(_gnd_net_),
            .in3(N__47612),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_16_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_16_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_16_20_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43118),
            .in3(N__46825),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53771),
            .ce(),
            .sr(N__53366));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47613),
            .lcout(\current_shift_inst.N_1619_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_20_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_20_6  (
            .in0(N__47615),
            .in1(N__46529),
            .in2(_gnd_net_),
            .in3(N__43295),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_20_7 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_20_7  (
            .in0(N__46502),
            .in1(N__47616),
            .in2(_gnd_net_),
            .in3(N__43283),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_16_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_16_21_0 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_16_21_0  (
            .in0(N__46919),
            .in1(N__47665),
            .in2(_gnd_net_),
            .in3(N__43274),
            .lcout(\current_shift_inst.control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_21_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_21_1  (
            .in0(N__47664),
            .in1(N__46583),
            .in2(_gnd_net_),
            .in3(N__43262),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_16_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_16_21_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_16_21_2  (
            .in0(N__47651),
            .in1(N__46964),
            .in2(_gnd_net_),
            .in3(N__43253),
            .lcout(\current_shift_inst.control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_3  (
            .in0(N__46661),
            .in1(N__43244),
            .in2(_gnd_net_),
            .in3(N__47649),
            .lcout(\current_shift_inst.control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_16_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_16_21_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_16_21_4  (
            .in0(N__47652),
            .in1(N__43235),
            .in2(_gnd_net_),
            .in3(N__46868),
            .lcout(\current_shift_inst.control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_21_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_21_5  (
            .in0(N__46733),
            .in1(N__43223),
            .in2(_gnd_net_),
            .in3(N__47648),
            .lcout(\current_shift_inst.control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_21_6 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_21_6  (
            .in0(N__47647),
            .in1(_gnd_net_),
            .in2(N__43211),
            .in3(N__46775),
            .lcout(\current_shift_inst.control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_21_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_21_7  (
            .in0(N__43199),
            .in1(N__46634),
            .in2(_gnd_net_),
            .in3(N__47650),
            .lcout(\current_shift_inst.control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_16_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_16_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43435),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53760),
            .ce(),
            .sr(N__53375));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_16_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_16_22_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_16_22_6  (
            .in0(N__52236),
            .in1(N__47858),
            .in2(_gnd_net_),
            .in3(N__52421),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53760),
            .ce(),
            .sr(N__53375));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_16_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_16_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43411),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53760),
            .ce(),
            .sr(N__53375));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_16_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_16_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47698),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_16_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_16_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_16_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_16_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43381),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53749),
            .ce(),
            .sr(N__53387));
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_16_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_16_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_16_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_28_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43360),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53749),
            .ce(),
            .sr(N__53387));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_16_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_16_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_16_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43339),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53749),
            .ce(),
            .sr(N__53387));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_16_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_16_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_16_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43309),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53749),
            .ce(),
            .sr(N__53387));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_16_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_16_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_16_24_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_16_24_5  (
            .in0(N__52420),
            .in1(N__47897),
            .in2(_gnd_net_),
            .in3(N__52238),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53749),
            .ce(),
            .sr(N__53387));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_16_24_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_16_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_16_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_16_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43519),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53749),
            .ce(),
            .sr(N__53387));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_16_24_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_16_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_16_24_7 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_16_24_7  (
            .in0(N__52419),
            .in1(N__47918),
            .in2(_gnd_net_),
            .in3(N__52237),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53749),
            .ce(),
            .sr(N__53387));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_16_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_16_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_16_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_16_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43495),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53744),
            .ce(),
            .sr(N__53393));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_16_25_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_16_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_16_25_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_16_25_1  (
            .in0(N__52368),
            .in1(N__48047),
            .in2(_gnd_net_),
            .in3(N__52215),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53744),
            .ce(),
            .sr(N__53393));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_16_25_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_16_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_16_25_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_16_25_2  (
            .in0(N__43462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53744),
            .ce(),
            .sr(N__53393));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_25_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_25_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_16_25_3  (
            .in0(N__52371),
            .in1(N__52214),
            .in2(_gnd_net_),
            .in3(N__48263),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53744),
            .ce(),
            .sr(N__53393));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_25_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_16_25_4  (
            .in0(N__52211),
            .in1(N__52373),
            .in2(_gnd_net_),
            .in3(N__48239),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53744),
            .ce(),
            .sr(N__53393));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_25_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_25_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_16_25_5  (
            .in0(N__52369),
            .in1(N__52212),
            .in2(_gnd_net_),
            .in3(N__48377),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53744),
            .ce(),
            .sr(N__53393));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_25_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_16_25_6  (
            .in0(N__52210),
            .in1(N__52372),
            .in2(_gnd_net_),
            .in3(N__48290),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53744),
            .ce(),
            .sr(N__53393));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_16_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_16_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_16_25_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_16_25_7  (
            .in0(N__52370),
            .in1(N__52213),
            .in2(_gnd_net_),
            .in3(N__48317),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53744),
            .ce(),
            .sr(N__53393));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_26_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_26_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_16_26_0  (
            .in0(N__52204),
            .in1(N__52363),
            .in2(_gnd_net_),
            .in3(N__48557),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53740),
            .ce(),
            .sr(N__53404));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_26_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_26_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_16_26_2  (
            .in0(N__52206),
            .in1(N__52365),
            .in2(_gnd_net_),
            .in3(N__48485),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53740),
            .ce(),
            .sr(N__53404));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_26_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_26_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_16_26_3  (
            .in0(N__52362),
            .in1(N__52209),
            .in2(_gnd_net_),
            .in3(N__48512),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53740),
            .ce(),
            .sr(N__53404));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_26_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_26_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_26_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_16_26_4  (
            .in0(N__52207),
            .in1(N__52366),
            .in2(_gnd_net_),
            .in3(N__48461),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53740),
            .ce(),
            .sr(N__53404));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_26_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_26_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_16_26_5  (
            .in0(N__52361),
            .in1(N__52208),
            .in2(_gnd_net_),
            .in3(N__48215),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53740),
            .ce(),
            .sr(N__53404));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_16_26_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_16_26_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_16_26_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_16_26_6  (
            .in0(N__52205),
            .in1(N__52364),
            .in2(_gnd_net_),
            .in3(N__48536),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53740),
            .ce(),
            .sr(N__53404));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_16_27_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_16_27_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_16_27_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_16_27_2  (
            .in0(N__50950),
            .in1(N__51231),
            .in2(N__50848),
            .in3(N__50786),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_16_27_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_16_27_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_16_27_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_16_27_5  (
            .in0(N__51230),
            .in1(N__50840),
            .in2(N__50793),
            .in3(N__50949),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_16_27_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_16_27_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_16_27_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_16_27_6  (
            .in0(N__51140),
            .in1(N__51188),
            .in2(N__50681),
            .in3(N__51062),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_16_28_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_16_28_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_16_28_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_16_28_0  (
            .in0(N__52187),
            .in1(N__52401),
            .in2(_gnd_net_),
            .in3(N__48077),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53731),
            .ce(),
            .sr(N__53412));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_16_28_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_16_28_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_16_28_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_16_28_7  (
            .in0(N__52400),
            .in1(N__48104),
            .in2(_gnd_net_),
            .in3(N__52188),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53731),
            .ce(),
            .sr(N__53412));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_3_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_3_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_3_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_3_0  (
            .in0(_gnd_net_),
            .in1(N__44149),
            .in2(N__44093),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_17_3_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__53855),
            .ce(N__44194),
            .sr(N__53312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_3_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_3_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_3_1  (
            .in0(_gnd_net_),
            .in1(N__44545),
            .in2(N__44123),
            .in3(N__43658),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__53855),
            .ce(N__44194),
            .sr(N__53312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_3_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_3_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_3_2  (
            .in0(_gnd_net_),
            .in1(N__44092),
            .in2(N__44521),
            .in3(N__43637),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__53855),
            .ce(N__44194),
            .sr(N__53312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_3_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_3_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_3_3  (
            .in0(_gnd_net_),
            .in1(N__44546),
            .in2(N__44491),
            .in3(N__43616),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__53855),
            .ce(N__44194),
            .sr(N__53312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_3_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_3_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_3_4  (
            .in0(_gnd_net_),
            .in1(N__44458),
            .in2(N__44522),
            .in3(N__43586),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__53855),
            .ce(N__44194),
            .sr(N__53312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_3_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_3_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_3_5  (
            .in0(_gnd_net_),
            .in1(N__44428),
            .in2(N__44492),
            .in3(N__43559),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__53855),
            .ce(N__44194),
            .sr(N__53312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_3_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_3_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_3_6  (
            .in0(_gnd_net_),
            .in1(N__44395),
            .in2(N__44462),
            .in3(N__43529),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__53855),
            .ce(N__44194),
            .sr(N__53312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_3_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_3_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_3_7  (
            .in0(_gnd_net_),
            .in1(N__44362),
            .in2(N__44432),
            .in3(N__43868),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__53855),
            .ce(N__44194),
            .sr(N__53312));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_4_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_4_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_4_0  (
            .in0(_gnd_net_),
            .in1(N__44338),
            .in2(N__44402),
            .in3(N__43847),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_17_4_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__53854),
            .ce(N__44195),
            .sr(N__53313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_4_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_4_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_4_1  (
            .in0(_gnd_net_),
            .in1(N__44314),
            .in2(N__44369),
            .in3(N__43826),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__53854),
            .ce(N__44195),
            .sr(N__53313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_4_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_4_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_4_2  (
            .in0(_gnd_net_),
            .in1(N__44339),
            .in2(N__44776),
            .in3(N__43805),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__53854),
            .ce(N__44195),
            .sr(N__53313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_4_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_4_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_4_3  (
            .in0(_gnd_net_),
            .in1(N__44315),
            .in2(N__44746),
            .in3(N__43784),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__53854),
            .ce(N__44195),
            .sr(N__53313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_4_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_4_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_4_4  (
            .in0(_gnd_net_),
            .in1(N__44713),
            .in2(N__44777),
            .in3(N__43763),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__53854),
            .ce(N__44195),
            .sr(N__53313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_4_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_4_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_4_5  (
            .in0(_gnd_net_),
            .in1(N__44686),
            .in2(N__44747),
            .in3(N__43745),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__53854),
            .ce(N__44195),
            .sr(N__53313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_4_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_4_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_4_6  (
            .in0(_gnd_net_),
            .in1(N__44656),
            .in2(N__44717),
            .in3(N__43721),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__53854),
            .ce(N__44195),
            .sr(N__53313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_4_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_4_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_4_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_4_7  (
            .in0(_gnd_net_),
            .in1(N__44687),
            .in2(N__44626),
            .in3(N__43697),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__53854),
            .ce(N__44195),
            .sr(N__53313));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_5_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_5_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(N__44593),
            .in2(N__44663),
            .in3(N__44045),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_17_5_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__53853),
            .ce(N__44193),
            .sr(N__53315));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_5_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_5_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_5_1  (
            .in0(_gnd_net_),
            .in1(N__44569),
            .in2(N__44630),
            .in3(N__44024),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__53853),
            .ce(N__44193),
            .sr(N__53315));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_5_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_5_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_5_2  (
            .in0(_gnd_net_),
            .in1(N__44594),
            .in2(N__45013),
            .in3(N__44003),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__53853),
            .ce(N__44193),
            .sr(N__53315));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_5_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_5_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_5_3  (
            .in0(_gnd_net_),
            .in1(N__44570),
            .in2(N__44986),
            .in3(N__43982),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__53853),
            .ce(N__44193),
            .sr(N__53315));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_5_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_5_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_5_4  (
            .in0(_gnd_net_),
            .in1(N__44956),
            .in2(N__45014),
            .in3(N__43958),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__53853),
            .ce(N__44193),
            .sr(N__53315));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_5_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_5_5  (
            .in0(_gnd_net_),
            .in1(N__44929),
            .in2(N__44987),
            .in3(N__43937),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__53853),
            .ce(N__44193),
            .sr(N__53315));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_5_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_5_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_5_6  (
            .in0(_gnd_net_),
            .in1(N__44899),
            .in2(N__44960),
            .in3(N__43913),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__53853),
            .ce(N__44193),
            .sr(N__53315));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_5_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_5_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_5_7  (
            .in0(_gnd_net_),
            .in1(N__44866),
            .in2(N__44933),
            .in3(N__43892),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__53853),
            .ce(N__44193),
            .sr(N__53315));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_6_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_6_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__44839),
            .in2(N__44906),
            .in3(N__44273),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__53850),
            .ce(N__44182),
            .sr(N__53316));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_6_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_6_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(N__44818),
            .in2(N__44873),
            .in3(N__44252),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__53850),
            .ce(N__44182),
            .sr(N__53316));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_6_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(N__44840),
            .in2(N__44798),
            .in3(N__44237),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__53850),
            .ce(N__44182),
            .sr(N__53316));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_6_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_6_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_6_3  (
            .in0(_gnd_net_),
            .in1(N__44819),
            .in2(N__45287),
            .in3(N__44219),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__53850),
            .ce(N__44182),
            .sr(N__53316));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44216),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53850),
            .ce(N__44182),
            .sr(N__53316));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_7_0  (
            .in0(N__45395),
            .in1(N__44142),
            .in2(_gnd_net_),
            .in3(N__44126),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__53846),
            .ce(N__45268),
            .sr(N__53317));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_7_1  (
            .in0(N__45390),
            .in1(N__44115),
            .in2(_gnd_net_),
            .in3(N__44096),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__53846),
            .ce(N__45268),
            .sr(N__53317));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_7_2  (
            .in0(N__45396),
            .in1(N__44082),
            .in2(_gnd_net_),
            .in3(N__44066),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__53846),
            .ce(N__45268),
            .sr(N__53317));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_7_3  (
            .in0(N__45391),
            .in1(N__44539),
            .in2(_gnd_net_),
            .in3(N__44525),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__53846),
            .ce(N__45268),
            .sr(N__53317));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_7_4  (
            .in0(N__45397),
            .in1(N__44509),
            .in2(_gnd_net_),
            .in3(N__44495),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__53846),
            .ce(N__45268),
            .sr(N__53317));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_7_5  (
            .in0(N__45392),
            .in1(N__44479),
            .in2(_gnd_net_),
            .in3(N__44465),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__53846),
            .ce(N__45268),
            .sr(N__53317));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_7_6  (
            .in0(N__45394),
            .in1(N__44451),
            .in2(_gnd_net_),
            .in3(N__44435),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__53846),
            .ce(N__45268),
            .sr(N__53317));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_7_7  (
            .in0(N__45393),
            .in1(N__44421),
            .in2(_gnd_net_),
            .in3(N__44405),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__53846),
            .ce(N__45268),
            .sr(N__53317));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_8_0  (
            .in0(N__45381),
            .in1(N__44394),
            .in2(_gnd_net_),
            .in3(N__44372),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__53841),
            .ce(N__45251),
            .sr(N__53318));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_8_1  (
            .in0(N__45407),
            .in1(N__44361),
            .in2(_gnd_net_),
            .in3(N__44342),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__53841),
            .ce(N__45251),
            .sr(N__53318));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_8_2  (
            .in0(N__45378),
            .in1(N__44332),
            .in2(_gnd_net_),
            .in3(N__44318),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__53841),
            .ce(N__45251),
            .sr(N__53318));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_8_3  (
            .in0(N__45404),
            .in1(N__44308),
            .in2(_gnd_net_),
            .in3(N__44294),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__53841),
            .ce(N__45251),
            .sr(N__53318));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_8_4  (
            .in0(N__45379),
            .in1(N__44764),
            .in2(_gnd_net_),
            .in3(N__44750),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__53841),
            .ce(N__45251),
            .sr(N__53318));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_8_5  (
            .in0(N__45405),
            .in1(N__44734),
            .in2(_gnd_net_),
            .in3(N__44720),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__53841),
            .ce(N__45251),
            .sr(N__53318));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_8_6  (
            .in0(N__45380),
            .in1(N__44706),
            .in2(_gnd_net_),
            .in3(N__44690),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__53841),
            .ce(N__45251),
            .sr(N__53318));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_8_7  (
            .in0(N__45406),
            .in1(N__44680),
            .in2(_gnd_net_),
            .in3(N__44666),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__53841),
            .ce(N__45251),
            .sr(N__53318));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_9_0  (
            .in0(N__45382),
            .in1(N__44655),
            .in2(_gnd_net_),
            .in3(N__44633),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__53834),
            .ce(N__45269),
            .sr(N__53320));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_9_1  (
            .in0(N__45386),
            .in1(N__44619),
            .in2(_gnd_net_),
            .in3(N__44597),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__53834),
            .ce(N__45269),
            .sr(N__53320));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_9_2  (
            .in0(N__45383),
            .in1(N__44587),
            .in2(_gnd_net_),
            .in3(N__44573),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__53834),
            .ce(N__45269),
            .sr(N__53320));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_9_3  (
            .in0(N__45387),
            .in1(N__44563),
            .in2(_gnd_net_),
            .in3(N__44549),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__53834),
            .ce(N__45269),
            .sr(N__53320));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_9_4  (
            .in0(N__45384),
            .in1(N__45006),
            .in2(_gnd_net_),
            .in3(N__44990),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__53834),
            .ce(N__45269),
            .sr(N__53320));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_9_5  (
            .in0(N__45388),
            .in1(N__44979),
            .in2(_gnd_net_),
            .in3(N__44963),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__53834),
            .ce(N__45269),
            .sr(N__53320));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_9_6  (
            .in0(N__45385),
            .in1(N__44955),
            .in2(_gnd_net_),
            .in3(N__44936),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__53834),
            .ce(N__45269),
            .sr(N__53320));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_9_7  (
            .in0(N__45389),
            .in1(N__44928),
            .in2(_gnd_net_),
            .in3(N__44909),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__53834),
            .ce(N__45269),
            .sr(N__53320));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_10_0  (
            .in0(N__45398),
            .in1(N__44898),
            .in2(_gnd_net_),
            .in3(N__44876),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__53829),
            .ce(N__45267),
            .sr(N__53322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_10_1  (
            .in0(N__45402),
            .in1(N__44865),
            .in2(_gnd_net_),
            .in3(N__44843),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__53829),
            .ce(N__45267),
            .sr(N__53322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_10_2  (
            .in0(N__45399),
            .in1(N__44838),
            .in2(_gnd_net_),
            .in3(N__44822),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__53829),
            .ce(N__45267),
            .sr(N__53322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_10_3  (
            .in0(N__45403),
            .in1(N__44817),
            .in2(_gnd_net_),
            .in3(N__44801),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__53829),
            .ce(N__45267),
            .sr(N__53322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_10_4  (
            .in0(N__45400),
            .in1(N__44794),
            .in2(_gnd_net_),
            .in3(N__44780),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__53829),
            .ce(N__45267),
            .sr(N__53322));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_10_5  (
            .in0(N__45283),
            .in1(N__45401),
            .in2(_gnd_net_),
            .in3(N__45290),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53829),
            .ce(N__45267),
            .sr(N__53322));
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_17_11_0  (
            .in0(N__48769),
            .in1(N__45216),
            .in2(_gnd_net_),
            .in3(N__45194),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__53823),
            .ce(N__48824),
            .sr(N__53324));
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_17_11_1  (
            .in0(N__48765),
            .in1(N__45180),
            .in2(_gnd_net_),
            .in3(N__45155),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__53823),
            .ce(N__48824),
            .sr(N__53324));
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_17_11_2  (
            .in0(N__48770),
            .in1(N__45145),
            .in2(_gnd_net_),
            .in3(N__45131),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__53823),
            .ce(N__48824),
            .sr(N__53324));
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_17_11_3  (
            .in0(N__48766),
            .in1(N__45121),
            .in2(_gnd_net_),
            .in3(N__45107),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__53823),
            .ce(N__48824),
            .sr(N__53324));
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_17_11_4  (
            .in0(N__48771),
            .in1(N__45091),
            .in2(_gnd_net_),
            .in3(N__45077),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__53823),
            .ce(N__48824),
            .sr(N__53324));
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_17_11_5  (
            .in0(N__48767),
            .in1(N__45061),
            .in2(_gnd_net_),
            .in3(N__45047),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__53823),
            .ce(N__48824),
            .sr(N__53324));
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_17_11_6  (
            .in0(N__48772),
            .in1(N__45033),
            .in2(_gnd_net_),
            .in3(N__45017),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__53823),
            .ce(N__48824),
            .sr(N__53324));
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_17_11_7  (
            .in0(N__48768),
            .in1(N__45637),
            .in2(_gnd_net_),
            .in3(N__45623),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__53823),
            .ce(N__48824),
            .sr(N__53324));
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_17_12_0  (
            .in0(N__48751),
            .in1(N__45615),
            .in2(_gnd_net_),
            .in3(N__45587),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__53815),
            .ce(N__48816),
            .sr(N__53328));
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_17_12_1  (
            .in0(N__48776),
            .in1(N__45570),
            .in2(_gnd_net_),
            .in3(N__45548),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__53815),
            .ce(N__48816),
            .sr(N__53328));
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_17_12_2  (
            .in0(N__48748),
            .in1(N__45534),
            .in2(_gnd_net_),
            .in3(N__45518),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__53815),
            .ce(N__48816),
            .sr(N__53328));
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_17_12_3  (
            .in0(N__48773),
            .in1(N__45508),
            .in2(_gnd_net_),
            .in3(N__45494),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__53815),
            .ce(N__48816),
            .sr(N__53328));
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_17_12_4  (
            .in0(N__48749),
            .in1(N__45484),
            .in2(_gnd_net_),
            .in3(N__45470),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__53815),
            .ce(N__48816),
            .sr(N__53328));
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_17_12_5  (
            .in0(N__48774),
            .in1(N__45454),
            .in2(_gnd_net_),
            .in3(N__45440),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__53815),
            .ce(N__48816),
            .sr(N__53328));
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_17_12_6  (
            .in0(N__48750),
            .in1(N__45424),
            .in2(_gnd_net_),
            .in3(N__45410),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__53815),
            .ce(N__48816),
            .sr(N__53328));
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_17_12_7  (
            .in0(N__48775),
            .in1(N__45904),
            .in2(_gnd_net_),
            .in3(N__45890),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__53815),
            .ce(N__48816),
            .sr(N__53328));
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_17_13_0  (
            .in0(N__48744),
            .in1(N__45882),
            .in2(_gnd_net_),
            .in3(N__45854),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__53807),
            .ce(N__48815),
            .sr(N__53330));
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_17_13_1  (
            .in0(N__48752),
            .in1(N__45843),
            .in2(_gnd_net_),
            .in3(N__45815),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__53807),
            .ce(N__48815),
            .sr(N__53330));
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_17_13_2  (
            .in0(N__48745),
            .in1(N__45801),
            .in2(_gnd_net_),
            .in3(N__45785),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__53807),
            .ce(N__48815),
            .sr(N__53330));
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_17_13_3  (
            .in0(N__48753),
            .in1(N__45775),
            .in2(_gnd_net_),
            .in3(N__45761),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__53807),
            .ce(N__48815),
            .sr(N__53330));
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_17_13_4  (
            .in0(N__48746),
            .in1(N__45747),
            .in2(_gnd_net_),
            .in3(N__45731),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__53807),
            .ce(N__48815),
            .sr(N__53330));
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_17_13_5  (
            .in0(N__48754),
            .in1(N__45715),
            .in2(_gnd_net_),
            .in3(N__45701),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__53807),
            .ce(N__48815),
            .sr(N__53330));
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_17_13_6  (
            .in0(N__48747),
            .in1(N__45687),
            .in2(_gnd_net_),
            .in3(N__45671),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__53807),
            .ce(N__48815),
            .sr(N__53330));
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_17_13_7  (
            .in0(N__48755),
            .in1(N__45661),
            .in2(_gnd_net_),
            .in3(N__45647),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__53807),
            .ce(N__48815),
            .sr(N__53330));
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_17_14_0  (
            .in0(N__48720),
            .in1(N__46158),
            .in2(_gnd_net_),
            .in3(N__46136),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__53800),
            .ce(N__48817),
            .sr(N__53336));
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_17_14_1  (
            .in0(N__48724),
            .in1(N__46125),
            .in2(_gnd_net_),
            .in3(N__46097),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__53800),
            .ce(N__48817),
            .sr(N__53336));
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_17_14_2  (
            .in0(N__48721),
            .in1(N__46087),
            .in2(_gnd_net_),
            .in3(N__46073),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__53800),
            .ce(N__48817),
            .sr(N__53336));
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_17_14_3  (
            .in0(N__48725),
            .in1(N__46063),
            .in2(_gnd_net_),
            .in3(N__46049),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__53800),
            .ce(N__48817),
            .sr(N__53336));
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_17_14_4  (
            .in0(N__48722),
            .in1(N__46036),
            .in2(_gnd_net_),
            .in3(N__46022),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__53800),
            .ce(N__48817),
            .sr(N__53336));
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_17_14_5  (
            .in0(N__46009),
            .in1(N__48723),
            .in2(_gnd_net_),
            .in3(N__46019),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53800),
            .ce(N__48817),
            .sr(N__53336));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__45995),
            .in2(N__45979),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__45930),
            .in2(N__45959),
            .in3(N__46425),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_15_2  (
            .in0(N__46426),
            .in1(N__49314),
            .in2(N__46376),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__50171),
            .in2(N__49499),
            .in3(N__46346),
            .lcout(\current_shift_inst.un38_control_input_0_s0_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__49318),
            .in2(N__46343),
            .in3(N__46316),
            .lcout(\current_shift_inst.un38_control_input_0_s0_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__46313),
            .in2(N__49500),
            .in3(N__46289),
            .lcout(\current_shift_inst.un38_control_input_0_s0_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__49322),
            .in2(N__46286),
            .in3(N__46259),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__46256),
            .in2(N__49501),
            .in3(N__46232),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__49342),
            .in2(N__46229),
            .in3(N__46199),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__46196),
            .in2(N__49506),
            .in3(N__46172),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__49346),
            .in2(N__46619),
            .in3(N__46595),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__46592),
            .in2(N__49507),
            .in3(N__46571),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__49350),
            .in2(N__46568),
            .in3(N__46544),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__46541),
            .in2(N__49508),
            .in3(N__46517),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__49354),
            .in2(N__46514),
            .in3(N__46490),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__46487),
            .in2(N__49509),
            .in3(N__46469),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__49510),
            .in2(N__46466),
            .in3(N__46442),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__46439),
            .in2(N__49615),
            .in3(N__46793),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__49514),
            .in2(N__46790),
            .in3(N__46763),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__46760),
            .in2(N__49616),
            .in3(N__46748),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__49518),
            .in2(N__46745),
            .in3(N__46718),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__46715),
            .in2(N__49617),
            .in3(N__46700),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__49522),
            .in2(N__46697),
            .in3(N__46676),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__46673),
            .in2(N__49618),
            .in3(N__46649),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__49526),
            .in2(N__46646),
            .in3(N__46622),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__46997),
            .in2(N__49619),
            .in3(N__46979),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__49530),
            .in2(N__46976),
            .in3(N__46952),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__46949),
            .in2(N__49620),
            .in3(N__46937),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__49534),
            .in2(N__46934),
            .in3(N__46910),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__46907),
            .in2(N__49621),
            .in3(N__46886),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(N__49538),
            .in2(N__46883),
            .in3(N__46859),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_18_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_18_7  (
            .in0(N__46856),
            .in1(N__46844),
            .in2(N__47687),
            .in3(N__46835),
            .lcout(\current_shift_inst.control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_17_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_17_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__46832),
            .in2(N__46826),
            .in3(N__46824),
            .lcout(\current_shift_inst.control_input_1 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_17_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_17_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__47165),
            .in2(_gnd_net_),
            .in3(N__47147),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_17_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_17_19_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__47144),
            .in2(_gnd_net_),
            .in3(N__47126),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_17_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_17_19_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__47123),
            .in2(_gnd_net_),
            .in3(N__47105),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_17_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_17_19_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__47102),
            .in2(_gnd_net_),
            .in3(N__47084),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_17_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_17_19_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__47081),
            .in2(_gnd_net_),
            .in3(N__47063),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_17_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_17_19_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__47060),
            .in2(_gnd_net_),
            .in3(N__47042),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_17_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_17_19_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(N__47039),
            .in2(_gnd_net_),
            .in3(N__47021),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_17_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_17_20_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__47018),
            .in2(_gnd_net_),
            .in3(N__47000),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_17_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_17_20_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__47345),
            .in2(_gnd_net_),
            .in3(N__47327),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_17_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_17_20_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__47324),
            .in2(_gnd_net_),
            .in3(N__47306),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_17_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_17_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__47303),
            .in2(_gnd_net_),
            .in3(N__47285),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_17_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_17_20_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__47282),
            .in2(_gnd_net_),
            .in3(N__47261),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_17_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_17_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__47258),
            .in2(_gnd_net_),
            .in3(N__47237),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_12 ),
            .carryout(\current_shift_inst.control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_17_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_17_20_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__47234),
            .in2(_gnd_net_),
            .in3(N__47213),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_13 ),
            .carryout(\current_shift_inst.control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_17_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_17_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__47210),
            .in2(_gnd_net_),
            .in3(N__47192),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_14 ),
            .carryout(\current_shift_inst.control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_17_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_17_21_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(N__47189),
            .in2(_gnd_net_),
            .in3(N__47168),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\current_shift_inst.control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_17_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_17_21_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__47519),
            .in2(_gnd_net_),
            .in3(N__47501),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_16 ),
            .carryout(\current_shift_inst.control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_17_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_17_21_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__47498),
            .in2(_gnd_net_),
            .in3(N__47474),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_17 ),
            .carryout(\current_shift_inst.control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_17_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_17_21_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(N__47471),
            .in2(_gnd_net_),
            .in3(N__47447),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_18 ),
            .carryout(\current_shift_inst.control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_17_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_17_21_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(N__47444),
            .in2(_gnd_net_),
            .in3(N__47426),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_19 ),
            .carryout(\current_shift_inst.control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_17_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_17_21_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(N__47423),
            .in2(_gnd_net_),
            .in3(N__47405),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_20 ),
            .carryout(\current_shift_inst.control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_17_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_17_21_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(N__47402),
            .in2(_gnd_net_),
            .in3(N__47381),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_21 ),
            .carryout(\current_shift_inst.control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_17_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_17_21_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(N__47378),
            .in2(_gnd_net_),
            .in3(N__47360),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_22 ),
            .carryout(\current_shift_inst.control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_17_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_17_22_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(N__47357),
            .in2(_gnd_net_),
            .in3(N__47819),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(\current_shift_inst.control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_17_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_17_22_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_17_22_1  (
            .in0(_gnd_net_),
            .in1(N__47816),
            .in2(_gnd_net_),
            .in3(N__47798),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_24 ),
            .carryout(\current_shift_inst.control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_17_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_17_22_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(N__47795),
            .in2(_gnd_net_),
            .in3(N__47771),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_25 ),
            .carryout(\current_shift_inst.control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_17_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_17_22_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(N__47768),
            .in2(_gnd_net_),
            .in3(N__47750),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_26 ),
            .carryout(\current_shift_inst.control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_17_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_17_22_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_17_22_4  (
            .in0(_gnd_net_),
            .in1(N__47747),
            .in2(_gnd_net_),
            .in3(N__47726),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_27 ),
            .carryout(\current_shift_inst.control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_17_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_17_22_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(N__47543),
            .in2(_gnd_net_),
            .in3(N__47711),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_28 ),
            .carryout(\current_shift_inst.control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_17_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_17_22_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_17_22_6  (
            .in0(N__47686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47708),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_17_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_17_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_17_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47685),
            .lcout(\current_shift_inst.control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_17_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_17_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_17_23_0 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_17_23_0  (
            .in0(_gnd_net_),
            .in1(N__51518),
            .in2(N__47537),
            .in3(N__52223),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(N__53761),
            .ce(),
            .sr(N__53376));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_17_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_17_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_17_23_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_17_23_1  (
            .in0(N__52222),
            .in1(N__51555),
            .in2(N__47996),
            .in3(N__47978),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(N__53761),
            .ce(),
            .sr(N__53376));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_17_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_17_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_17_23_2 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_17_23_2  (
            .in0(N__52235),
            .in1(N__51618),
            .in2(N__47975),
            .in3(N__47957),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(N__53761),
            .ce(),
            .sr(N__53376));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(N__51595),
            .in2(N__47954),
            .in3(N__47936),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(N__51771),
            .in2(N__47933),
            .in3(N__47912),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(N__51804),
            .in2(N__47909),
            .in3(N__47891),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(N__51315),
            .in2(N__47888),
            .in3(N__47873),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_23_7  (
            .in0(_gnd_net_),
            .in1(N__51474),
            .in2(N__47870),
            .in3(N__47852),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_24_0  (
            .in0(_gnd_net_),
            .in1(N__47849),
            .in2(N__51280),
            .in3(N__47834),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__50749),
            .in2(N__48206),
            .in3(N__48176),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_24_2  (
            .in0(_gnd_net_),
            .in1(N__51378),
            .in2(N__48173),
            .in3(N__48155),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_24_3  (
            .in0(_gnd_net_),
            .in1(N__50685),
            .in2(N__48152),
            .in3(N__48122),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_24_4  (
            .in0(_gnd_net_),
            .in1(N__50629),
            .in2(N__48119),
            .in3(N__48092),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_24_5  (
            .in0(_gnd_net_),
            .in1(N__50578),
            .in2(N__48089),
            .in3(N__48065),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_24_6  (
            .in0(_gnd_net_),
            .in1(N__50522),
            .in2(N__48062),
            .in3(N__48041),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(N__52068),
            .in2(N__48038),
            .in3(N__48020),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_25_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_25_0  (
            .in0(_gnd_net_),
            .in1(N__52462),
            .in2(N__48017),
            .in3(N__47999),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_17_25_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_25_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_25_1  (
            .in0(_gnd_net_),
            .in1(N__51436),
            .in2(N__48416),
            .in3(N__48398),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_25_2  (
            .in0(_gnd_net_),
            .in1(N__51689),
            .in2(N__48395),
            .in3(N__48371),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_25_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_25_3  (
            .in0(_gnd_net_),
            .in1(N__51748),
            .in2(N__48368),
            .in3(N__48338),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_25_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_25_4  (
            .in0(_gnd_net_),
            .in1(N__50945),
            .in2(N__48335),
            .in3(N__48311),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_25_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_25_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_25_5  (
            .in0(_gnd_net_),
            .in1(N__51656),
            .in2(N__48308),
            .in3(N__48284),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_25_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_25_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_25_6  (
            .in0(_gnd_net_),
            .in1(N__50905),
            .in2(N__48281),
            .in3(N__48257),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_25_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_25_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_25_7  (
            .in0(_gnd_net_),
            .in1(N__48254),
            .in2(N__50844),
            .in3(N__48233),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_26_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_26_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_26_0  (
            .in0(_gnd_net_),
            .in1(N__48230),
            .in2(N__50794),
            .in3(N__48209),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_17_26_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_26_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_26_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_26_1  (
            .in0(_gnd_net_),
            .in1(N__51232),
            .in2(N__48575),
            .in3(N__48551),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_26_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_26_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_26_2  (
            .in0(_gnd_net_),
            .in1(N__48548),
            .in2(N__51196),
            .in3(N__48530),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_26_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_26_3  (
            .in0(_gnd_net_),
            .in1(N__48527),
            .in2(N__51148),
            .in3(N__48506),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_26_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_26_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_26_4  (
            .in0(_gnd_net_),
            .in1(N__51096),
            .in2(N__48503),
            .in3(N__48479),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_26_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_26_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_26_5  (
            .in0(_gnd_net_),
            .in1(N__48476),
            .in2(N__51070),
            .in3(N__48455),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_17_26_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_17_26_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_17_26_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_er_31_LC_17_26_6  (
            .in0(N__52374),
            .in1(N__48452),
            .in2(N__48437),
            .in3(N__48419),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53745),
            .ce(N__52221),
            .sr(N__53394));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_17_27_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_17_27_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_17_27_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_17_27_0  (
            .in0(N__50904),
            .in1(N__50526),
            .in2(N__51100),
            .in3(N__50747),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_17_27_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_17_27_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_17_27_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_17_27_1  (
            .in0(N__51746),
            .in1(N__51660),
            .in2(N__51707),
            .in3(N__52454),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_17_27_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_17_27_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_17_27_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_17_27_2  (
            .in0(N__51379),
            .in1(N__50571),
            .in2(N__52073),
            .in3(N__50622),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_17_27_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_17_27_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_17_27_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_17_27_3  (
            .in0(N__48650),
            .in1(N__48644),
            .in2(N__48638),
            .in3(N__48635),
            .lcout(\current_shift_inst.PI_CTRL.N_46_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_17_27_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_17_27_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_17_27_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_17_27_4  (
            .in0(N__51063),
            .in1(N__51141),
            .in2(N__50692),
            .in3(N__51189),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_17_27_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_17_27_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_17_27_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_17_27_5  (
            .in0(_gnd_net_),
            .in1(N__51092),
            .in2(_gnd_net_),
            .in3(N__50903),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_17_27_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_17_27_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_17_27_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_17_27_6  (
            .in0(N__48629),
            .in1(N__50527),
            .in2(N__48620),
            .in3(N__50748),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_17_28_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_17_28_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_17_28_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_17_28_2  (
            .in0(N__48617),
            .in1(N__52388),
            .in2(_gnd_net_),
            .in3(N__52189),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53733),
            .ce(),
            .sr(N__53408));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_17_28_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_17_28_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_17_28_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_17_28_3  (
            .in0(N__51432),
            .in1(N__48884),
            .in2(N__52418),
            .in3(N__48608),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_17_28_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_17_28_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_17_28_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_17_28_4  (
            .in0(N__48602),
            .in1(N__48593),
            .in2(N__48587),
            .in3(N__51449),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_17_28_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_17_28_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_17_28_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_17_28_5  (
            .in0(N__51008),
            .in1(N__51401),
            .in2(N__48584),
            .in3(N__48581),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_17_28_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_17_28_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_17_28_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_17_28_6  (
            .in0(_gnd_net_),
            .in1(N__52387),
            .in2(N__48899),
            .in3(N__48896),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53733),
            .ce(),
            .sr(N__53408));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_17_29_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_17_29_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_17_29_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_17_29_4  (
            .in0(N__50570),
            .in1(N__50618),
            .in2(N__51377),
            .in3(N__52058),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_18_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_18_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48870),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48833),
            .ce(),
            .sr(N__53325));
    defparam \delay_measurement_inst.stop_timer_tr_LC_18_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_18_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_18_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48871),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48833),
            .ce(),
            .sr(N__53325));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_13_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_13_3  (
            .in0(N__48791),
            .in1(N__49062),
            .in2(_gnd_net_),
            .in3(N__49031),
            .lcout(\current_shift_inst.timer_s1.N_164_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_18_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_18_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_18_14_2 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_18_14_2  (
            .in0(N__49084),
            .in1(N__49144),
            .in2(N__49037),
            .in3(N__48793),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53808),
            .ce(),
            .sr(N__53331));
    defparam \current_shift_inst.timer_s1.running_LC_18_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_18_14_3 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_18_14_3  (
            .in0(N__48794),
            .in1(N__49032),
            .in2(_gnd_net_),
            .in3(N__49063),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53808),
            .ce(),
            .sr(N__53331));
    defparam \current_shift_inst.start_timer_s1_LC_18_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_18_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_18_14_6 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_18_14_6  (
            .in0(N__49083),
            .in1(N__48792),
            .in2(_gnd_net_),
            .in3(N__49145),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53808),
            .ce(),
            .sr(N__53331));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49061),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_18_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_18_15_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_18_15_6  (
            .in0(N__50082),
            .in1(N__49804),
            .in2(N__49562),
            .in3(N__50164),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_15_7 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_15_7  (
            .in0(N__50165),
            .in1(N__50081),
            .in2(N__49805),
            .in3(N__49459),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S1_LC_18_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_18_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_18_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49143),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53793),
            .ce(),
            .sr(N__53338));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_18_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_18_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__49064),
            .in2(_gnd_net_),
            .in3(N__49036),
            .lcout(\current_shift_inst.timer_s1.N_163_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_18_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_18_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__50185),
            .in2(_gnd_net_),
            .in3(N__51534),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53781),
            .ce(),
            .sr(N__53355));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_18_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_18_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_18_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48982),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53776),
            .ce(),
            .sr(N__53362));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_18_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_18_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_18_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48964),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53776),
            .ce(),
            .sr(N__53362));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_18_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_18_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_18_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_18_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48940),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53776),
            .ce(),
            .sr(N__53362));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_18_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_18_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_18_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_18_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48919),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53776),
            .ce(),
            .sr(N__53362));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_18_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_18_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_18_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50374),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53772),
            .ce(),
            .sr(N__53367));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_18_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_18_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_18_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50353),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53772),
            .ce(),
            .sr(N__53367));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_18_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_18_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_18_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50329),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53772),
            .ce(),
            .sr(N__53367));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_18_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_18_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_18_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50302),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53772),
            .ce(),
            .sr(N__53367));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_18_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_18_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_18_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_18_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50278),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53772),
            .ce(),
            .sr(N__53367));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_18_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_18_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_18_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_18_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50257),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53772),
            .ce(),
            .sr(N__53367));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_18_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_18_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_18_22_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_18_22_6  (
            .in0(N__50233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53772),
            .ce(),
            .sr(N__53367));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_18_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_18_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_18_22_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_18_22_7  (
            .in0(N__50206),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53772),
            .ce(),
            .sr(N__53367));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_18_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_18_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_18_23_0  (
            .in0(_gnd_net_),
            .in1(N__50186),
            .in2(N__51535),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_23_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_18_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_18_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_18_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(N__50468),
            .in2(N__51562),
            .in3(N__50462),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__53765),
            .ce(),
            .sr(N__53370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_18_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_18_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_18_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_18_23_2  (
            .in0(_gnd_net_),
            .in1(N__51622),
            .in2(N__50459),
            .in3(N__50450),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__53765),
            .ce(),
            .sr(N__53370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_18_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_18_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_18_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(N__50447),
            .in2(N__51602),
            .in3(N__50438),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__53765),
            .ce(),
            .sr(N__53370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_18_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_18_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_18_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__50435),
            .in2(N__51785),
            .in3(N__50423),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__53765),
            .ce(),
            .sr(N__53370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_18_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_18_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_18_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_18_23_5  (
            .in0(_gnd_net_),
            .in1(N__50420),
            .in2(N__51818),
            .in3(N__50411),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__53765),
            .ce(),
            .sr(N__53370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_18_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_18_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_18_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(N__50408),
            .in2(N__51332),
            .in3(N__50399),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__53765),
            .ce(),
            .sr(N__53370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_18_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_18_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_18_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(N__50396),
            .in2(N__51500),
            .in3(N__50390),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__53765),
            .ce(),
            .sr(N__53370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_18_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_18_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_18_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_18_24_0  (
            .in0(_gnd_net_),
            .in1(N__50387),
            .in2(N__51281),
            .in3(N__50378),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_18_24_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__53762),
            .ce(),
            .sr(N__53377));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_18_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_18_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_18_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_18_24_1  (
            .in0(_gnd_net_),
            .in1(N__50762),
            .in2(N__50753),
            .in3(N__50720),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__53762),
            .ce(),
            .sr(N__53377));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_18_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_18_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_18_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_18_24_2  (
            .in0(_gnd_net_),
            .in1(N__50717),
            .in2(N__51383),
            .in3(N__50708),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__53762),
            .ce(),
            .sr(N__53377));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_18_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_18_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_18_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_18_24_3  (
            .in0(_gnd_net_),
            .in1(N__50705),
            .in2(N__50696),
            .in3(N__50648),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__53762),
            .ce(),
            .sr(N__53377));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_18_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_18_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_18_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_18_24_4  (
            .in0(_gnd_net_),
            .in1(N__50645),
            .in2(N__50636),
            .in3(N__50594),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__53762),
            .ce(),
            .sr(N__53377));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_18_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_18_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_18_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_18_24_5  (
            .in0(_gnd_net_),
            .in1(N__50591),
            .in2(N__50582),
            .in3(N__50549),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__53762),
            .ce(),
            .sr(N__53377));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_18_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_18_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_18_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_18_24_6  (
            .in0(_gnd_net_),
            .in1(N__50546),
            .in2(N__50534),
            .in3(N__50501),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__53762),
            .ce(),
            .sr(N__53377));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_18_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_18_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_18_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_18_24_7  (
            .in0(_gnd_net_),
            .in1(N__50498),
            .in2(N__52072),
            .in3(N__50489),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__53762),
            .ce(),
            .sr(N__53377));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_18_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_18_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_18_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_18_25_0  (
            .in0(_gnd_net_),
            .in1(N__50486),
            .in2(N__52466),
            .in3(N__50471),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_18_25_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__53754),
            .ce(),
            .sr(N__53383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_18_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_18_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_18_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_18_25_1  (
            .in0(_gnd_net_),
            .in1(N__51002),
            .in2(N__51443),
            .in3(N__50993),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__53754),
            .ce(),
            .sr(N__53383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_18_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_18_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_18_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_18_25_2  (
            .in0(_gnd_net_),
            .in1(N__50990),
            .in2(N__51706),
            .in3(N__50978),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__53754),
            .ce(),
            .sr(N__53383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_18_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_18_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_18_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_18_25_3  (
            .in0(_gnd_net_),
            .in1(N__50975),
            .in2(N__51752),
            .in3(N__50966),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__53754),
            .ce(),
            .sr(N__53383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_18_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_18_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_18_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_18_25_4  (
            .in0(_gnd_net_),
            .in1(N__50963),
            .in2(N__50954),
            .in3(N__50924),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__53754),
            .ce(),
            .sr(N__53383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_18_25_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_18_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_18_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_18_25_5  (
            .in0(_gnd_net_),
            .in1(N__51664),
            .in2(N__50921),
            .in3(N__50909),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__53754),
            .ce(),
            .sr(N__53383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_18_25_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_18_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_18_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_18_25_6  (
            .in0(_gnd_net_),
            .in1(N__50906),
            .in2(N__50879),
            .in3(N__50864),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__53754),
            .ce(),
            .sr(N__53383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_18_25_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_18_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_18_25_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_18_25_7  (
            .in0(_gnd_net_),
            .in1(N__50861),
            .in2(N__50849),
            .in3(N__50813),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__53754),
            .ce(),
            .sr(N__53383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_18_26_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_18_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_18_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_18_26_0  (
            .in0(_gnd_net_),
            .in1(N__50810),
            .in2(N__50801),
            .in3(N__50765),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_18_26_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__53750),
            .ce(),
            .sr(N__53388));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_18_26_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_18_26_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_18_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_18_26_1  (
            .in0(_gnd_net_),
            .in1(N__51248),
            .in2(N__51239),
            .in3(N__51212),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__53750),
            .ce(),
            .sr(N__53388));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_18_26_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_18_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_18_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_18_26_2  (
            .in0(_gnd_net_),
            .in1(N__51209),
            .in2(N__51200),
            .in3(N__51167),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__53750),
            .ce(),
            .sr(N__53388));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_18_26_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_18_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_18_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_18_26_3  (
            .in0(_gnd_net_),
            .in1(N__51164),
            .in2(N__51152),
            .in3(N__51119),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__53750),
            .ce(),
            .sr(N__53388));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_18_26_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_18_26_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_18_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_18_26_4  (
            .in0(_gnd_net_),
            .in1(N__51116),
            .in2(N__51104),
            .in3(N__51074),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__53750),
            .ce(),
            .sr(N__53388));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_18_26_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_18_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_18_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_18_26_5  (
            .in0(_gnd_net_),
            .in1(N__51071),
            .in2(N__51041),
            .in3(N__51026),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__53750),
            .ce(),
            .sr(N__53388));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_18_26_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_18_26_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_18_26_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_18_26_6  (
            .in0(N__52367),
            .in1(N__51023),
            .in2(_gnd_net_),
            .in3(N__51014),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53750),
            .ce(),
            .sr(N__53388));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_18_27_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_18_27_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_18_27_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_18_27_0  (
            .in0(N__51275),
            .in1(N__51814),
            .in2(N__51331),
            .in3(N__51781),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_18_27_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_18_27_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_18_27_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_18_27_1  (
            .in0(N__51629),
            .in1(N__51496),
            .in2(N__51011),
            .in3(N__51594),
            .lcout(\current_shift_inst.PI_CTRL.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_18_27_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_18_27_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_18_27_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_18_27_2  (
            .in0(N__51324),
            .in1(N__51813),
            .in2(_gnd_net_),
            .in3(N__51780),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_18_27_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_18_27_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_18_27_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_18_27_4  (
            .in0(N__51747),
            .in1(N__51705),
            .in2(N__51668),
            .in3(N__52455),
            .lcout(\current_shift_inst.PI_CTRL.N_46_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_18_27_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_18_27_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_18_27_5 .LUT_INIT=16'b0001000100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_18_27_5  (
            .in0(N__51628),
            .in1(N__51593),
            .in2(N__51569),
            .in3(N__51539),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_18_27_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_18_27_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_18_27_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_18_27_6  (
            .in0(N__51276),
            .in1(N__51495),
            .in2(N__51458),
            .in3(N__51455),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_18_28_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_18_28_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_18_28_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_18_28_0  (
            .in0(N__52375),
            .in1(N__51431),
            .in2(_gnd_net_),
            .in3(N__51407),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_18_29_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_18_29_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_18_29_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_18_29_6  (
            .in0(N__52422),
            .in1(N__51395),
            .in2(_gnd_net_),
            .in3(N__52190),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53734),
            .ce(),
            .sr(N__53409));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_20_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_20_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_20_23_3 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_20_23_3  (
            .in0(N__52425),
            .in1(N__51341),
            .in2(_gnd_net_),
            .in3(N__52234),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53777),
            .ce(),
            .sr(N__53371));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_20_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_20_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_20_23_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_20_23_4  (
            .in0(N__52233),
            .in1(N__52426),
            .in2(_gnd_net_),
            .in3(N__51293),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53777),
            .ce(),
            .sr(N__53371));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_20_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_20_24_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_20_24_0  (
            .in0(_gnd_net_),
            .in1(N__51877),
            .in2(_gnd_net_),
            .in3(N__51859),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_20_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_20_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_20_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_20_24_1  (
            .in0(N__52009),
            .in1(N__52022),
            .in2(N__51989),
            .in3(N__51974),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_20_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_20_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_20_24_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_20_24_2  (
            .in0(N__52021),
            .in1(N__51928),
            .in2(N__52010),
            .in3(N__51949),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_20_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_20_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_20_24_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_20_24_3  (
            .in0(N__51985),
            .in1(N__51973),
            .in2(N__51962),
            .in3(N__51959),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_20_25_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_20_25_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_20_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_20_25_0  (
            .in0(N__52622),
            .in1(N__51953),
            .in2(N__51935),
            .in3(N__52601),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_20_25_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_20_25_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_20_25_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_20_25_2  (
            .in0(N__51907),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52648),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_20_25_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_20_25_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_20_25_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_20_25_3  (
            .in0(N__51896),
            .in1(N__51842),
            .in2(N__51911),
            .in3(N__51830),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_20_25_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_20_25_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_20_25_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_20_25_4  (
            .in0(N__51908),
            .in1(N__51895),
            .in2(N__51884),
            .in3(N__51863),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_20_25_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_20_25_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_20_25_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_20_25_5  (
            .in0(_gnd_net_),
            .in1(N__51841),
            .in2(_gnd_net_),
            .in3(N__51829),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_20_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_20_25_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_20_25_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_20_25_6  (
            .in0(N__52579),
            .in1(N__52658),
            .in2(N__52652),
            .in3(N__52649),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_20_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_20_25_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_20_25_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_20_25_7  (
            .in0(N__52637),
            .in1(N__52631),
            .in2(N__52625),
            .in3(N__52484),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_20_26_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_20_26_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_20_26_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_20_26_0  (
            .in0(N__52531),
            .in1(N__52519),
            .in2(N__52505),
            .in3(N__52621),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_20_26_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_20_26_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_20_26_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_20_26_4  (
            .in0(N__52544),
            .in1(N__52600),
            .in2(N__52559),
            .in3(N__52580),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_20_26_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_20_26_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_20_26_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_20_26_5  (
            .in0(_gnd_net_),
            .in1(N__52558),
            .in2(_gnd_net_),
            .in3(N__52543),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_20_26_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_20_26_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_20_26_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_20_26_6  (
            .in0(N__52532),
            .in1(N__52520),
            .in2(N__52508),
            .in3(N__52504),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_20_27_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_20_27_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_20_27_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_20_27_6  (
            .in0(N__52424),
            .in1(N__52478),
            .in2(_gnd_net_),
            .in3(N__52241),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53755),
            .ce(),
            .sr(N__53395));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_21_25_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_21_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_21_25_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_21_25_1  (
            .in0(N__52427),
            .in1(N__52253),
            .in2(_gnd_net_),
            .in3(N__52239),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53773),
            .ce(),
            .sr(N__53389));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_22_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_22_25_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_22_25_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_22_25_7  (
            .in0(N__52901),
            .in1(N__52889),
            .in2(N__52880),
            .in3(N__52865),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_23_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_23_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_23_15_5 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_23_15_5  (
            .in0(N__54085),
            .in1(N__53993),
            .in2(N__52838),
            .in3(N__54259),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53835),
            .ce(),
            .sr(N__53343));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_23_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_23_17_3 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_23_17_3  (
            .in0(N__52831),
            .in1(N__53002),
            .in2(N__53056),
            .in3(N__52802),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(\current_shift_inst.PI_CTRL.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_17_4 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_23_17_4  (
            .in0(N__54063),
            .in1(N__54165),
            .in2(N__52841),
            .in3(N__54246),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_18_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_23_18_0  (
            .in0(_gnd_net_),
            .in1(N__52830),
            .in2(_gnd_net_),
            .in3(N__53043),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_18_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_23_18_1  (
            .in0(N__52989),
            .in1(N__52699),
            .in2(N__52805),
            .in3(N__53093),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_23_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_23_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_23_18_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_23_18_5  (
            .in0(_gnd_net_),
            .in1(N__52698),
            .in2(_gnd_net_),
            .in3(N__53092),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_0  (
            .in0(N__54091),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_duty_input_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53842),
            .ce(),
            .sr(N__53347));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_15_3 .LUT_INIT=16'b1000100011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_24_15_3  (
            .in0(N__52703),
            .in1(N__53992),
            .in2(N__54260),
            .in3(N__54092),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53842),
            .ce(),
            .sr(N__53347));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_16_0 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_24_16_0  (
            .in0(N__54261),
            .in1(N__54089),
            .in2(N__53994),
            .in3(N__53091),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53836),
            .ce(),
            .sr(N__53356));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_1 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_1  (
            .in0(N__54088),
            .in1(N__53982),
            .in2(N__53057),
            .in3(N__54263),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53836),
            .ce(),
            .sr(N__53356));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_16_2 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_24_16_2  (
            .in0(N__54262),
            .in1(N__54090),
            .in2(N__53995),
            .in3(N__53003),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53836),
            .ce(),
            .sr(N__53356));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_3 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_3  (
            .in0(N__54116),
            .in1(N__53915),
            .in2(_gnd_net_),
            .in3(N__54191),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53836),
            .ce(),
            .sr(N__53356));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4  (
            .in0(_gnd_net_),
            .in1(N__53900),
            .in2(_gnd_net_),
            .in3(N__54177),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53836),
            .ce(),
            .sr(N__53356));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_5 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_5  (
            .in0(N__52907),
            .in1(N__54167),
            .in2(N__53996),
            .in3(N__54014),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53836),
            .ce(),
            .sr(N__53356));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_24_16_6  (
            .in0(_gnd_net_),
            .in1(N__52946),
            .in2(_gnd_net_),
            .in3(N__54178),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53836),
            .ce(),
            .sr(N__53356));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_24_16_7  (
            .in0(N__54179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52928),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53836),
            .ce(),
            .sr(N__53356));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_24_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_24_17_3 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_24_17_3  (
            .in0(N__54166),
            .in1(N__54087),
            .in2(N__54278),
            .in3(N__54248),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_24_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_24_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_24_17_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_24_17_5  (
            .in0(N__54274),
            .in1(N__54086),
            .in2(_gnd_net_),
            .in3(N__54247),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_17_6 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_24_17_6  (
            .in0(N__54115),
            .in1(N__53911),
            .in2(N__54194),
            .in3(N__54190),
            .lcout(\current_shift_inst.PI_CTRL.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_24_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_24_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_24_18_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_24_18_4  (
            .in0(_gnd_net_),
            .in1(N__54164),
            .in2(_gnd_net_),
            .in3(N__54114),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_18_5 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_24_18_5  (
            .in0(N__54067),
            .in1(N__54010),
            .in2(N__53999),
            .in3(N__53965),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_24_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53861),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53816),
            .ce(),
            .sr(N__53372));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_24_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_24_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_24_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_24_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53890),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53816),
            .ce(),
            .sr(N__53372));
endmodule // MAIN
